../sin_cos.sv