module ghost (
    input   [11:0]  address,
    input     clock,
    output reg [11:0]  q
);

reg [11:0]mem[0:((1 << $bits(address))-1)];
reg [11:0]address_q;

initial
begin
	mem[12'h000] = 12'hFFF;
	mem[12'h001] = 12'hFFF;
	mem[12'h002] = 12'hFFF;
	mem[12'h003] = 12'hFFF;
	mem[12'h004] = 12'hFFF;
	mem[12'h005] = 12'hFFF;
	mem[12'h006] = 12'hFFF;
	mem[12'h007] = 12'hFFF;
	mem[12'h008] = 12'hFFF;
	mem[12'h009] = 12'hFFF;
	mem[12'h00A] = 12'hFFF;
	mem[12'h00B] = 12'hFFF;
	mem[12'h00C] = 12'hFFF;
	mem[12'h00D] = 12'hFFF;
	mem[12'h00E] = 12'hFFF;
	mem[12'h00F] = 12'hFFF;
	mem[12'h010] = 12'hFFF;
	mem[12'h011] = 12'hFFF;
	mem[12'h012] = 12'hFFF;
	mem[12'h013] = 12'hFFF;
	mem[12'h014] = 12'hFFF;
	mem[12'h015] = 12'hFFF;
	mem[12'h016] = 12'hFFF;
	mem[12'h017] = 12'hFFF;
	mem[12'h018] = 12'hFFF;
	mem[12'h019] = 12'hFFF;
	mem[12'h01A] = 12'hFFF;
	mem[12'h01B] = 12'hFFF;
	mem[12'h01C] = 12'hFFF;
	mem[12'h01D] = 12'hFFF;
	mem[12'h01E] = 12'hFFF;
	mem[12'h01F] = 12'hFFF;
	mem[12'h020] = 12'hFFF;
	mem[12'h021] = 12'hFFF;
	mem[12'h022] = 12'hFFF;
	mem[12'h023] = 12'hFFF;
	mem[12'h024] = 12'hFFF;
	mem[12'h025] = 12'hFFF;
	mem[12'h026] = 12'hFFF;
	mem[12'h027] = 12'hFFF;
	mem[12'h028] = 12'hFFF;
	mem[12'h029] = 12'hFFF;
	mem[12'h02A] = 12'hFFF;
	mem[12'h02B] = 12'hFFF;
	mem[12'h02C] = 12'hFFF;
	mem[12'h02D] = 12'hFFF;
	mem[12'h02E] = 12'hFFF;
	mem[12'h02F] = 12'hFFF;
	mem[12'h030] = 12'hFFF;
	mem[12'h031] = 12'hFFF;
	mem[12'h032] = 12'hFFF;
	mem[12'h033] = 12'hFFF;
	mem[12'h034] = 12'hFFF;
	mem[12'h035] = 12'hFFF;
	mem[12'h036] = 12'hFFF;
	mem[12'h037] = 12'hFFF;
	mem[12'h038] = 12'hFFF;
	mem[12'h039] = 12'hFFF;
	mem[12'h03A] = 12'hFFF;
	mem[12'h03B] = 12'hFFF;
	mem[12'h03C] = 12'hFFF;
	mem[12'h03D] = 12'hFFF;
	mem[12'h03E] = 12'hFFF;
	mem[12'h03F] = 12'hFFF;
	mem[12'h040] = 12'hFFF;
	mem[12'h041] = 12'hFFF;
	mem[12'h042] = 12'hFFF;
	mem[12'h043] = 12'hFFF;
	mem[12'h044] = 12'hFFF;
	mem[12'h045] = 12'hFFF;
	mem[12'h046] = 12'hFFF;
	mem[12'h047] = 12'hFFF;
	mem[12'h048] = 12'hFFF;
	mem[12'h049] = 12'hFFF;
	mem[12'h04A] = 12'hFFF;
	mem[12'h04B] = 12'hFFF;
	mem[12'h04C] = 12'hFFF;
	mem[12'h04D] = 12'hFFF;
	mem[12'h04E] = 12'hFFF;
	mem[12'h04F] = 12'hFFF;
	mem[12'h050] = 12'hFFF;
	mem[12'h051] = 12'hFFF;
	mem[12'h052] = 12'hFFF;
	mem[12'h053] = 12'hFFF;
	mem[12'h054] = 12'hFFF;
	mem[12'h055] = 12'hFFF;
	mem[12'h056] = 12'hFFF;
	mem[12'h057] = 12'hFFF;
	mem[12'h058] = 12'hFFF;
	mem[12'h059] = 12'hFFF;
	mem[12'h05A] = 12'hFFF;
	mem[12'h05B] = 12'hFFF;
	mem[12'h05C] = 12'hFFF;
	mem[12'h05D] = 12'hFFF;
	mem[12'h05E] = 12'hFFF;
	mem[12'h05F] = 12'hFFF;
	mem[12'h060] = 12'hFFF;
	mem[12'h061] = 12'hFFF;
	mem[12'h062] = 12'hFFF;
	mem[12'h063] = 12'hFFF;
	mem[12'h064] = 12'hFFF;
	mem[12'h065] = 12'hFFF;
	mem[12'h066] = 12'hFFF;
	mem[12'h067] = 12'hFFF;
	mem[12'h068] = 12'hFFF;
	mem[12'h069] = 12'hFFF;
	mem[12'h06A] = 12'hFFF;
	mem[12'h06B] = 12'hFFF;
	mem[12'h06C] = 12'hFFF;
	mem[12'h06D] = 12'hFFF;
	mem[12'h06E] = 12'hFFF;
	mem[12'h06F] = 12'hFFF;
	mem[12'h070] = 12'hFFF;
	mem[12'h071] = 12'hFFF;
	mem[12'h072] = 12'hFFF;
	mem[12'h073] = 12'hFFF;
	mem[12'h074] = 12'hFFF;
	mem[12'h075] = 12'hFFF;
	mem[12'h076] = 12'hFFF;
	mem[12'h077] = 12'hFFF;
	mem[12'h078] = 12'hFFF;
	mem[12'h079] = 12'hFFF;
	mem[12'h07A] = 12'hFFF;
	mem[12'h07B] = 12'hFFF;
	mem[12'h07C] = 12'hFFF;
	mem[12'h07D] = 12'hFFF;
	mem[12'h07E] = 12'hFFF;
	mem[12'h07F] = 12'hFFF;
	mem[12'h080] = 12'hFFF;
	mem[12'h081] = 12'hFFF;
	mem[12'h082] = 12'hFFF;
	mem[12'h083] = 12'hFFF;
	mem[12'h084] = 12'hFFF;
	mem[12'h085] = 12'hFFF;
	mem[12'h086] = 12'hFFF;
	mem[12'h087] = 12'hFFF;
	mem[12'h088] = 12'hFFF;
	mem[12'h089] = 12'hFFF;
	mem[12'h08A] = 12'hFFF;
	mem[12'h08B] = 12'hFFF;
	mem[12'h08C] = 12'hFFF;
	mem[12'h08D] = 12'hFFF;
	mem[12'h08E] = 12'hFFF;
	mem[12'h08F] = 12'hFFF;
	mem[12'h090] = 12'hFFF;
	mem[12'h091] = 12'hFFF;
	mem[12'h092] = 12'hFFF;
	mem[12'h093] = 12'hFFF;
	mem[12'h094] = 12'hFFF;
	mem[12'h095] = 12'hFFF;
	mem[12'h096] = 12'hFFF;
	mem[12'h097] = 12'hFFF;
	mem[12'h098] = 12'hFFF;
	mem[12'h099] = 12'hFFF;
	mem[12'h09A] = 12'hFFF;
	mem[12'h09B] = 12'hFFF;
	mem[12'h09C] = 12'hFFF;
	mem[12'h09D] = 12'hFFF;
	mem[12'h09E] = 12'hFFF;
	mem[12'h09F] = 12'hFFF;
	mem[12'h0A0] = 12'hFFF;
	mem[12'h0A1] = 12'hFFF;
	mem[12'h0A2] = 12'hFFF;
	mem[12'h0A3] = 12'hFFF;
	mem[12'h0A4] = 12'hFFF;
	mem[12'h0A5] = 12'hFFF;
	mem[12'h0A6] = 12'hFFF;
	mem[12'h0A7] = 12'hFFF;
	mem[12'h0A8] = 12'hFFF;
	mem[12'h0A9] = 12'hFFF;
	mem[12'h0AA] = 12'hFFF;
	mem[12'h0AB] = 12'hFFF;
	mem[12'h0AC] = 12'hFFF;
	mem[12'h0AD] = 12'hFFF;
	mem[12'h0AE] = 12'hFFF;
	mem[12'h0AF] = 12'hFFF;
	mem[12'h0B0] = 12'hFFF;
	mem[12'h0B1] = 12'hFFF;
	mem[12'h0B2] = 12'hFFF;
	mem[12'h0B3] = 12'hFFF;
	mem[12'h0B4] = 12'hFFF;
	mem[12'h0B5] = 12'hFFF;
	mem[12'h0B6] = 12'hFFF;
	mem[12'h0B7] = 12'hFFF;
	mem[12'h0B8] = 12'hFFF;
	mem[12'h0B9] = 12'hFFF;
	mem[12'h0BA] = 12'hFFF;
	mem[12'h0BB] = 12'hFFF;
	mem[12'h0BC] = 12'hFFF;
	mem[12'h0BD] = 12'hFFF;
	mem[12'h0BE] = 12'hFFF;
	mem[12'h0BF] = 12'hFFF;
	mem[12'h0C0] = 12'hFFF;
	mem[12'h0C1] = 12'hFFF;
	mem[12'h0C2] = 12'hFFF;
	mem[12'h0C3] = 12'hFFF;
	mem[12'h0C4] = 12'hFFF;
	mem[12'h0C5] = 12'hFFF;
	mem[12'h0C6] = 12'hFFF;
	mem[12'h0C7] = 12'hFFF;
	mem[12'h0C8] = 12'hFFF;
	mem[12'h0C9] = 12'hFFF;
	mem[12'h0CA] = 12'hFFF;
	mem[12'h0CB] = 12'hFFF;
	mem[12'h0CC] = 12'hFFF;
	mem[12'h0CD] = 12'hFFF;
	mem[12'h0CE] = 12'hFFF;
	mem[12'h0CF] = 12'hFFF;
	mem[12'h0D0] = 12'hFFF;
	mem[12'h0D1] = 12'hFFF;
	mem[12'h0D2] = 12'hFFF;
	mem[12'h0D3] = 12'hFFF;
	mem[12'h0D4] = 12'hFFF;
	mem[12'h0D5] = 12'hFFF;
	mem[12'h0D6] = 12'hFFF;
	mem[12'h0D7] = 12'hFFF;
	mem[12'h0D8] = 12'hFFF;
	mem[12'h0D9] = 12'hFFF;
	mem[12'h0DA] = 12'hFFF;
	mem[12'h0DB] = 12'hFFF;
	mem[12'h0DC] = 12'hFFF;
	mem[12'h0DD] = 12'hFFF;
	mem[12'h0DE] = 12'hFFF;
	mem[12'h0DF] = 12'hFFF;
	mem[12'h0E0] = 12'hFFF;
	mem[12'h0E1] = 12'hFFF;
	mem[12'h0E2] = 12'hFFF;
	mem[12'h0E3] = 12'hFFF;
	mem[12'h0E4] = 12'hFFF;
	mem[12'h0E5] = 12'hFFF;
	mem[12'h0E6] = 12'hFFF;
	mem[12'h0E7] = 12'hFFF;
	mem[12'h0E8] = 12'hFFF;
	mem[12'h0E9] = 12'hFFF;
	mem[12'h0EA] = 12'hFFF;
	mem[12'h0EB] = 12'hFFF;
	mem[12'h0EC] = 12'hFFF;
	mem[12'h0ED] = 12'hFFF;
	mem[12'h0EE] = 12'hFFF;
	mem[12'h0EF] = 12'hFFF;
	mem[12'h0F0] = 12'hFFF;
	mem[12'h0F1] = 12'hFFF;
	mem[12'h0F2] = 12'hFFF;
	mem[12'h0F3] = 12'hFFF;
	mem[12'h0F4] = 12'hFFF;
	mem[12'h0F5] = 12'hFFF;
	mem[12'h0F6] = 12'hFFF;
	mem[12'h0F7] = 12'hFFF;
	mem[12'h0F8] = 12'hFFF;
	mem[12'h0F9] = 12'hFFF;
	mem[12'h0FA] = 12'hFFF;
	mem[12'h0FB] = 12'hFFF;
	mem[12'h0FC] = 12'hFFF;
	mem[12'h0FD] = 12'hFFF;
	mem[12'h0FE] = 12'hFFF;
	mem[12'h0FF] = 12'hFFF;
	mem[12'h100] = 12'hFFF;
	mem[12'h101] = 12'hFFF;
	mem[12'h102] = 12'hFFF;
	mem[12'h103] = 12'hFFF;
	mem[12'h104] = 12'hFFF;
	mem[12'h105] = 12'hFFF;
	mem[12'h106] = 12'hFFF;
	mem[12'h107] = 12'hFFF;
	mem[12'h108] = 12'hFFF;
	mem[12'h109] = 12'hFFF;
	mem[12'h10A] = 12'hFFF;
	mem[12'h10B] = 12'hFFF;
	mem[12'h10C] = 12'hFFF;
	mem[12'h10D] = 12'hFFF;
	mem[12'h10E] = 12'hFFF;
	mem[12'h10F] = 12'hFFF;
	mem[12'h110] = 12'hFFF;
	mem[12'h111] = 12'hFFF;
	mem[12'h112] = 12'hFFF;
	mem[12'h113] = 12'hFFF;
	mem[12'h114] = 12'hFFF;
	mem[12'h115] = 12'hFFF;
	mem[12'h116] = 12'hFFF;
	mem[12'h117] = 12'hFFF;
	mem[12'h118] = 12'hFFF;
	mem[12'h119] = 12'hFFF;
	mem[12'h11A] = 12'hFFF;
	mem[12'h11B] = 12'hF00;
	mem[12'h11C] = 12'hF00;
	mem[12'h11D] = 12'hF00;
	mem[12'h11E] = 12'hF00;
	mem[12'h11F] = 12'hF00;
	mem[12'h120] = 12'hF00;
	mem[12'h121] = 12'hF00;
	mem[12'h122] = 12'hF00;
	mem[12'h123] = 12'hF00;
	mem[12'h124] = 12'hF00;
	mem[12'h125] = 12'hFFF;
	mem[12'h126] = 12'hFFF;
	mem[12'h127] = 12'hFFF;
	mem[12'h128] = 12'hFFF;
	mem[12'h129] = 12'hFFF;
	mem[12'h12A] = 12'hFFF;
	mem[12'h12B] = 12'hFFF;
	mem[12'h12C] = 12'hFFF;
	mem[12'h12D] = 12'hFFF;
	mem[12'h12E] = 12'hFFF;
	mem[12'h12F] = 12'hFFF;
	mem[12'h130] = 12'hFFF;
	mem[12'h131] = 12'hFFF;
	mem[12'h132] = 12'hFFF;
	mem[12'h133] = 12'hFFF;
	mem[12'h134] = 12'hFFF;
	mem[12'h135] = 12'hFFF;
	mem[12'h136] = 12'hFFF;
	mem[12'h137] = 12'hFFF;
	mem[12'h138] = 12'hFFF;
	mem[12'h139] = 12'hFFF;
	mem[12'h13A] = 12'hFFF;
	mem[12'h13B] = 12'hFFF;
	mem[12'h13C] = 12'hFFF;
	mem[12'h13D] = 12'hFFF;
	mem[12'h13E] = 12'hFFF;
	mem[12'h13F] = 12'hFFF;
	mem[12'h140] = 12'hFFF;
	mem[12'h141] = 12'hFFF;
	mem[12'h142] = 12'hFFF;
	mem[12'h143] = 12'hFFF;
	mem[12'h144] = 12'hFFF;
	mem[12'h145] = 12'hFFF;
	mem[12'h146] = 12'hFFF;
	mem[12'h147] = 12'hFFF;
	mem[12'h148] = 12'hFFF;
	mem[12'h149] = 12'hFFF;
	mem[12'h14A] = 12'hFFF;
	mem[12'h14B] = 12'hFFF;
	mem[12'h14C] = 12'hFFF;
	mem[12'h14D] = 12'hFFF;
	mem[12'h14E] = 12'hFFF;
	mem[12'h14F] = 12'hFFF;
	mem[12'h150] = 12'hFFF;
	mem[12'h151] = 12'hFFF;
	mem[12'h152] = 12'hFFF;
	mem[12'h153] = 12'hFFF;
	mem[12'h154] = 12'hFFF;
	mem[12'h155] = 12'hFFF;
	mem[12'h156] = 12'hFFF;
	mem[12'h157] = 12'hFFF;
	mem[12'h158] = 12'hF00;
	mem[12'h159] = 12'hE22;
	mem[12'h15A] = 12'hE22;
	mem[12'h15B] = 12'hE22;
	mem[12'h15C] = 12'hF00;
	mem[12'h15D] = 12'hF00;
	mem[12'h15E] = 12'hF00;
	mem[12'h15F] = 12'hF00;
	mem[12'h160] = 12'hF00;
	mem[12'h161] = 12'hF00;
	mem[12'h162] = 12'hF00;
	mem[12'h163] = 12'hF00;
	mem[12'h164] = 12'hE22;
	mem[12'h165] = 12'hE22;
	mem[12'h166] = 12'hE22;
	mem[12'h167] = 12'hF00;
	mem[12'h168] = 12'hFFF;
	mem[12'h169] = 12'hFFF;
	mem[12'h16A] = 12'hFFF;
	mem[12'h16B] = 12'hFFF;
	mem[12'h16C] = 12'hFFF;
	mem[12'h16D] = 12'hFFF;
	mem[12'h16E] = 12'hFFF;
	mem[12'h16F] = 12'hFFF;
	mem[12'h170] = 12'hFFF;
	mem[12'h171] = 12'hFFF;
	mem[12'h172] = 12'hFFF;
	mem[12'h173] = 12'hFFF;
	mem[12'h174] = 12'hFFF;
	mem[12'h175] = 12'hFFF;
	mem[12'h176] = 12'hFFF;
	mem[12'h177] = 12'hFFF;
	mem[12'h178] = 12'hFFF;
	mem[12'h179] = 12'hFFF;
	mem[12'h17A] = 12'hFFF;
	mem[12'h17B] = 12'hFFF;
	mem[12'h17C] = 12'hFFF;
	mem[12'h17D] = 12'hFFF;
	mem[12'h17E] = 12'hFFF;
	mem[12'h17F] = 12'hFFF;
	mem[12'h180] = 12'hFFF;
	mem[12'h181] = 12'hFFF;
	mem[12'h182] = 12'hFFF;
	mem[12'h183] = 12'hFFF;
	mem[12'h184] = 12'hFFF;
	mem[12'h185] = 12'hFFF;
	mem[12'h186] = 12'hFFF;
	mem[12'h187] = 12'hFFF;
	mem[12'h188] = 12'hFFF;
	mem[12'h189] = 12'hFFF;
	mem[12'h18A] = 12'hFFF;
	mem[12'h18B] = 12'hFFF;
	mem[12'h18C] = 12'hFFF;
	mem[12'h18D] = 12'hFFF;
	mem[12'h18E] = 12'hFFF;
	mem[12'h18F] = 12'hFFF;
	mem[12'h190] = 12'hFFF;
	mem[12'h191] = 12'hFFF;
	mem[12'h192] = 12'hFFF;
	mem[12'h193] = 12'hFFF;
	mem[12'h194] = 12'hFFF;
	mem[12'h195] = 12'hF00;
	mem[12'h196] = 12'hE22;
	mem[12'h197] = 12'hE22;
	mem[12'h198] = 12'hF00;
	mem[12'h199] = 12'hF00;
	mem[12'h19A] = 12'hF00;
	mem[12'h19B] = 12'hF00;
	mem[12'h19C] = 12'hF00;
	mem[12'h19D] = 12'hF00;
	mem[12'h19E] = 12'hF00;
	mem[12'h19F] = 12'hF00;
	mem[12'h1A0] = 12'hF00;
	mem[12'h1A1] = 12'hF00;
	mem[12'h1A2] = 12'hF00;
	mem[12'h1A3] = 12'hF00;
	mem[12'h1A4] = 12'hF00;
	mem[12'h1A5] = 12'hF00;
	mem[12'h1A6] = 12'hF00;
	mem[12'h1A7] = 12'hF00;
	mem[12'h1A8] = 12'hE22;
	mem[12'h1A9] = 12'hE22;
	mem[12'h1AA] = 12'hF00;
	mem[12'h1AB] = 12'hFFF;
	mem[12'h1AC] = 12'hFFF;
	mem[12'h1AD] = 12'hFFF;
	mem[12'h1AE] = 12'hFFF;
	mem[12'h1AF] = 12'hFFF;
	mem[12'h1B0] = 12'hFFF;
	mem[12'h1B1] = 12'hFFF;
	mem[12'h1B2] = 12'hFFF;
	mem[12'h1B3] = 12'hFFF;
	mem[12'h1B4] = 12'hFFF;
	mem[12'h1B5] = 12'hFFF;
	mem[12'h1B6] = 12'hFFF;
	mem[12'h1B7] = 12'hFFF;
	mem[12'h1B8] = 12'hFFF;
	mem[12'h1B9] = 12'hFFF;
	mem[12'h1BA] = 12'hFFF;
	mem[12'h1BB] = 12'hFFF;
	mem[12'h1BC] = 12'hFFF;
	mem[12'h1BD] = 12'hFFF;
	mem[12'h1BE] = 12'hFFF;
	mem[12'h1BF] = 12'hFFF;
	mem[12'h1C0] = 12'hFFF;
	mem[12'h1C1] = 12'hFFF;
	mem[12'h1C2] = 12'hFFF;
	mem[12'h1C3] = 12'hFFF;
	mem[12'h1C4] = 12'hFFF;
	mem[12'h1C5] = 12'hFFF;
	mem[12'h1C6] = 12'hFFF;
	mem[12'h1C7] = 12'hFFF;
	mem[12'h1C8] = 12'hFFF;
	mem[12'h1C9] = 12'hFFF;
	mem[12'h1CA] = 12'hFFF;
	mem[12'h1CB] = 12'hFFF;
	mem[12'h1CC] = 12'hFFF;
	mem[12'h1CD] = 12'hFFF;
	mem[12'h1CE] = 12'hFFF;
	mem[12'h1CF] = 12'hFFF;
	mem[12'h1D0] = 12'hFFF;
	mem[12'h1D1] = 12'hFFF;
	mem[12'h1D2] = 12'hFFF;
	mem[12'h1D3] = 12'hF00;
	mem[12'h1D4] = 12'hE22;
	mem[12'h1D5] = 12'hE22;
	mem[12'h1D6] = 12'hF00;
	mem[12'h1D7] = 12'hF00;
	mem[12'h1D8] = 12'hF00;
	mem[12'h1D9] = 12'hF00;
	mem[12'h1DA] = 12'hF00;
	mem[12'h1DB] = 12'hF00;
	mem[12'h1DC] = 12'hF00;
	mem[12'h1DD] = 12'hF00;
	mem[12'h1DE] = 12'hF00;
	mem[12'h1DF] = 12'hF00;
	mem[12'h1E0] = 12'hF00;
	mem[12'h1E1] = 12'hF00;
	mem[12'h1E2] = 12'hF00;
	mem[12'h1E3] = 12'hF00;
	mem[12'h1E4] = 12'hF00;
	mem[12'h1E5] = 12'hF00;
	mem[12'h1E6] = 12'hF00;
	mem[12'h1E7] = 12'hF00;
	mem[12'h1E8] = 12'hF00;
	mem[12'h1E9] = 12'hF00;
	mem[12'h1EA] = 12'hE22;
	mem[12'h1EB] = 12'hE22;
	mem[12'h1EC] = 12'hF00;
	mem[12'h1ED] = 12'hFFF;
	mem[12'h1EE] = 12'hFFF;
	mem[12'h1EF] = 12'hFFF;
	mem[12'h1F0] = 12'hFFF;
	mem[12'h1F1] = 12'hFFF;
	mem[12'h1F2] = 12'hFFF;
	mem[12'h1F3] = 12'hFFF;
	mem[12'h1F4] = 12'hFFF;
	mem[12'h1F5] = 12'hFFF;
	mem[12'h1F6] = 12'hFFF;
	mem[12'h1F7] = 12'hFFF;
	mem[12'h1F8] = 12'hFFF;
	mem[12'h1F9] = 12'hFFF;
	mem[12'h1FA] = 12'hFFF;
	mem[12'h1FB] = 12'hFFF;
	mem[12'h1FC] = 12'hFFF;
	mem[12'h1FD] = 12'hFFF;
	mem[12'h1FE] = 12'hFFF;
	mem[12'h1FF] = 12'hFFF;
	mem[12'h200] = 12'hFFF;
	mem[12'h201] = 12'hFFF;
	mem[12'h202] = 12'hFFF;
	mem[12'h203] = 12'hFFF;
	mem[12'h204] = 12'hFFF;
	mem[12'h205] = 12'hFFF;
	mem[12'h206] = 12'hFFF;
	mem[12'h207] = 12'hFFF;
	mem[12'h208] = 12'hFFF;
	mem[12'h209] = 12'hFFF;
	mem[12'h20A] = 12'hFFF;
	mem[12'h20B] = 12'hFFF;
	mem[12'h20C] = 12'hFFF;
	mem[12'h20D] = 12'hFFF;
	mem[12'h20E] = 12'hFFF;
	mem[12'h20F] = 12'hFFF;
	mem[12'h210] = 12'hFFF;
	mem[12'h211] = 12'hE22;
	mem[12'h212] = 12'hE22;
	mem[12'h213] = 12'hF00;
	mem[12'h214] = 12'hF00;
	mem[12'h215] = 12'hF00;
	mem[12'h216] = 12'hF00;
	mem[12'h217] = 12'hF00;
	mem[12'h218] = 12'hF00;
	mem[12'h219] = 12'hF00;
	mem[12'h21A] = 12'hF00;
	mem[12'h21B] = 12'hF00;
	mem[12'h21C] = 12'hF00;
	mem[12'h21D] = 12'hF00;
	mem[12'h21E] = 12'hF00;
	mem[12'h21F] = 12'hF00;
	mem[12'h220] = 12'hF00;
	mem[12'h221] = 12'hF00;
	mem[12'h222] = 12'hF00;
	mem[12'h223] = 12'hF00;
	mem[12'h224] = 12'hF00;
	mem[12'h225] = 12'hF00;
	mem[12'h226] = 12'hF00;
	mem[12'h227] = 12'hF00;
	mem[12'h228] = 12'hF00;
	mem[12'h229] = 12'hF00;
	mem[12'h22A] = 12'hF00;
	mem[12'h22B] = 12'hF00;
	mem[12'h22C] = 12'hF00;
	mem[12'h22D] = 12'hE22;
	mem[12'h22E] = 12'hF00;
	mem[12'h22F] = 12'hFFF;
	mem[12'h230] = 12'hFFF;
	mem[12'h231] = 12'hFFF;
	mem[12'h232] = 12'hFFF;
	mem[12'h233] = 12'hFFF;
	mem[12'h234] = 12'hFFF;
	mem[12'h235] = 12'hFFF;
	mem[12'h236] = 12'hFFF;
	mem[12'h237] = 12'hFFF;
	mem[12'h238] = 12'hFFF;
	mem[12'h239] = 12'hFFF;
	mem[12'h23A] = 12'hFFF;
	mem[12'h23B] = 12'hFFF;
	mem[12'h23C] = 12'hFFF;
	mem[12'h23D] = 12'hFFF;
	mem[12'h23E] = 12'hFFF;
	mem[12'h23F] = 12'hFFF;
	mem[12'h240] = 12'hFFF;
	mem[12'h241] = 12'hFFF;
	mem[12'h242] = 12'hFFF;
	mem[12'h243] = 12'hFFF;
	mem[12'h244] = 12'hFFF;
	mem[12'h245] = 12'hFFF;
	mem[12'h246] = 12'hFFF;
	mem[12'h247] = 12'hFFF;
	mem[12'h248] = 12'hFFF;
	mem[12'h249] = 12'hFFF;
	mem[12'h24A] = 12'hFFF;
	mem[12'h24B] = 12'hFFF;
	mem[12'h24C] = 12'hFFF;
	mem[12'h24D] = 12'hFFF;
	mem[12'h24E] = 12'hFFF;
	mem[12'h24F] = 12'hFFF;
	mem[12'h250] = 12'hF00;
	mem[12'h251] = 12'hE22;
	mem[12'h252] = 12'hF00;
	mem[12'h253] = 12'hF00;
	mem[12'h254] = 12'hF00;
	mem[12'h255] = 12'hF00;
	mem[12'h256] = 12'hF00;
	mem[12'h257] = 12'hF00;
	mem[12'h258] = 12'hF00;
	mem[12'h259] = 12'hF00;
	mem[12'h25A] = 12'hF00;
	mem[12'h25B] = 12'hF00;
	mem[12'h25C] = 12'hF00;
	mem[12'h25D] = 12'hF00;
	mem[12'h25E] = 12'hF00;
	mem[12'h25F] = 12'hF00;
	mem[12'h260] = 12'hF00;
	mem[12'h261] = 12'hF00;
	mem[12'h262] = 12'hF00;
	mem[12'h263] = 12'hF00;
	mem[12'h264] = 12'hF00;
	mem[12'h265] = 12'hF00;
	mem[12'h266] = 12'hF00;
	mem[12'h267] = 12'hF00;
	mem[12'h268] = 12'hF00;
	mem[12'h269] = 12'hF00;
	mem[12'h26A] = 12'hF00;
	mem[12'h26B] = 12'hF00;
	mem[12'h26C] = 12'hF00;
	mem[12'h26D] = 12'hF00;
	mem[12'h26E] = 12'hE22;
	mem[12'h26F] = 12'hF00;
	mem[12'h270] = 12'hFFF;
	mem[12'h271] = 12'hFFF;
	mem[12'h272] = 12'hFFF;
	mem[12'h273] = 12'hFFF;
	mem[12'h274] = 12'hFFF;
	mem[12'h275] = 12'hFFF;
	mem[12'h276] = 12'hFFF;
	mem[12'h277] = 12'hFFF;
	mem[12'h278] = 12'hFFF;
	mem[12'h279] = 12'hFFF;
	mem[12'h27A] = 12'hFFF;
	mem[12'h27B] = 12'hFFF;
	mem[12'h27C] = 12'hFFF;
	mem[12'h27D] = 12'hFFF;
	mem[12'h27E] = 12'hFFF;
	mem[12'h27F] = 12'hFFF;
	mem[12'h280] = 12'hFFF;
	mem[12'h281] = 12'hFFF;
	mem[12'h282] = 12'hFFF;
	mem[12'h283] = 12'hFFF;
	mem[12'h284] = 12'hFFF;
	mem[12'h285] = 12'hFFF;
	mem[12'h286] = 12'hFFF;
	mem[12'h287] = 12'hFFF;
	mem[12'h288] = 12'hFFF;
	mem[12'h289] = 12'hFFF;
	mem[12'h28A] = 12'hFFF;
	mem[12'h28B] = 12'hFFF;
	mem[12'h28C] = 12'hFFF;
	mem[12'h28D] = 12'hFFF;
	mem[12'h28E] = 12'hFFF;
	mem[12'h28F] = 12'hF00;
	mem[12'h290] = 12'hF00;
	mem[12'h291] = 12'hF00;
	mem[12'h292] = 12'hF00;
	mem[12'h293] = 12'hF00;
	mem[12'h294] = 12'hF00;
	mem[12'h295] = 12'hF00;
	mem[12'h296] = 12'hF00;
	mem[12'h297] = 12'hF00;
	mem[12'h298] = 12'hF00;
	mem[12'h299] = 12'hF00;
	mem[12'h29A] = 12'hF00;
	mem[12'h29B] = 12'hF00;
	mem[12'h29C] = 12'hF00;
	mem[12'h29D] = 12'hF00;
	mem[12'h29E] = 12'hF00;
	mem[12'h29F] = 12'hF00;
	mem[12'h2A0] = 12'hF00;
	mem[12'h2A1] = 12'hF00;
	mem[12'h2A2] = 12'hF00;
	mem[12'h2A3] = 12'hF00;
	mem[12'h2A4] = 12'hF00;
	mem[12'h2A5] = 12'hF00;
	mem[12'h2A6] = 12'hF00;
	mem[12'h2A7] = 12'hF00;
	mem[12'h2A8] = 12'hF00;
	mem[12'h2A9] = 12'hF00;
	mem[12'h2AA] = 12'hF00;
	mem[12'h2AB] = 12'hF00;
	mem[12'h2AC] = 12'hF00;
	mem[12'h2AD] = 12'hF00;
	mem[12'h2AE] = 12'hF00;
	mem[12'h2AF] = 12'hF00;
	mem[12'h2B0] = 12'hF00;
	mem[12'h2B1] = 12'hFFF;
	mem[12'h2B2] = 12'hFFF;
	mem[12'h2B3] = 12'hFFF;
	mem[12'h2B4] = 12'hFFF;
	mem[12'h2B5] = 12'hFFF;
	mem[12'h2B6] = 12'hFFF;
	mem[12'h2B7] = 12'hFFF;
	mem[12'h2B8] = 12'hFFF;
	mem[12'h2B9] = 12'hFFF;
	mem[12'h2BA] = 12'hFFF;
	mem[12'h2BB] = 12'hFFF;
	mem[12'h2BC] = 12'hFFF;
	mem[12'h2BD] = 12'hFFF;
	mem[12'h2BE] = 12'hFFF;
	mem[12'h2BF] = 12'hFFF;
	mem[12'h2C0] = 12'hFFF;
	mem[12'h2C1] = 12'hFFF;
	mem[12'h2C2] = 12'hFFF;
	mem[12'h2C3] = 12'hFFF;
	mem[12'h2C4] = 12'hFFF;
	mem[12'h2C5] = 12'hFFF;
	mem[12'h2C6] = 12'hFFF;
	mem[12'h2C7] = 12'hFFF;
	mem[12'h2C8] = 12'hFFF;
	mem[12'h2C9] = 12'hFFF;
	mem[12'h2CA] = 12'hFFF;
	mem[12'h2CB] = 12'hFFF;
	mem[12'h2CC] = 12'hFFF;
	mem[12'h2CD] = 12'hFFF;
	mem[12'h2CE] = 12'hE22;
	mem[12'h2CF] = 12'hF00;
	mem[12'h2D0] = 12'hF00;
	mem[12'h2D1] = 12'hF00;
	mem[12'h2D2] = 12'hF00;
	mem[12'h2D3] = 12'hF00;
	mem[12'h2D4] = 12'hF00;
	mem[12'h2D5] = 12'hF00;
	mem[12'h2D6] = 12'hF00;
	mem[12'h2D7] = 12'hF00;
	mem[12'h2D8] = 12'hF00;
	mem[12'h2D9] = 12'hF00;
	mem[12'h2DA] = 12'hF00;
	mem[12'h2DB] = 12'hF00;
	mem[12'h2DC] = 12'hF00;
	mem[12'h2DD] = 12'hF00;
	mem[12'h2DE] = 12'hF00;
	mem[12'h2DF] = 12'hF00;
	mem[12'h2E0] = 12'hF00;
	mem[12'h2E1] = 12'hF00;
	mem[12'h2E2] = 12'hF00;
	mem[12'h2E3] = 12'hF00;
	mem[12'h2E4] = 12'hF00;
	mem[12'h2E5] = 12'hF00;
	mem[12'h2E6] = 12'hF00;
	mem[12'h2E7] = 12'hF00;
	mem[12'h2E8] = 12'hF00;
	mem[12'h2E9] = 12'hF00;
	mem[12'h2EA] = 12'hF00;
	mem[12'h2EB] = 12'hF00;
	mem[12'h2EC] = 12'hF00;
	mem[12'h2ED] = 12'hF00;
	mem[12'h2EE] = 12'hF00;
	mem[12'h2EF] = 12'hF00;
	mem[12'h2F0] = 12'hF00;
	mem[12'h2F1] = 12'hE22;
	mem[12'h2F2] = 12'hFFF;
	mem[12'h2F3] = 12'hFFF;
	mem[12'h2F4] = 12'hFFF;
	mem[12'h2F5] = 12'hFFF;
	mem[12'h2F6] = 12'hFFF;
	mem[12'h2F7] = 12'hFFF;
	mem[12'h2F8] = 12'hFFF;
	mem[12'h2F9] = 12'hFFF;
	mem[12'h2FA] = 12'hFFF;
	mem[12'h2FB] = 12'hFFF;
	mem[12'h2FC] = 12'hFFF;
	mem[12'h2FD] = 12'hFFF;
	mem[12'h2FE] = 12'hFFF;
	mem[12'h2FF] = 12'hFFF;
	mem[12'h300] = 12'hFFF;
	mem[12'h301] = 12'hFFF;
	mem[12'h302] = 12'hFFF;
	mem[12'h303] = 12'hFFF;
	mem[12'h304] = 12'hFFF;
	mem[12'h305] = 12'hFFF;
	mem[12'h306] = 12'hFFF;
	mem[12'h307] = 12'hFFF;
	mem[12'h308] = 12'hFFF;
	mem[12'h309] = 12'hFFF;
	mem[12'h30A] = 12'hFFF;
	mem[12'h30B] = 12'hFFF;
	mem[12'h30C] = 12'hFFF;
	mem[12'h30D] = 12'hF00;
	mem[12'h30E] = 12'hF00;
	mem[12'h30F] = 12'hF00;
	mem[12'h310] = 12'hF00;
	mem[12'h311] = 12'hF00;
	mem[12'h312] = 12'hF00;
	mem[12'h313] = 12'hF00;
	mem[12'h314] = 12'hF00;
	mem[12'h315] = 12'hF00;
	mem[12'h316] = 12'hF00;
	mem[12'h317] = 12'hF00;
	mem[12'h318] = 12'hF00;
	mem[12'h319] = 12'hF00;
	mem[12'h31A] = 12'hF00;
	mem[12'h31B] = 12'hF00;
	mem[12'h31C] = 12'hF00;
	mem[12'h31D] = 12'hF00;
	mem[12'h31E] = 12'hF00;
	mem[12'h31F] = 12'hF00;
	mem[12'h320] = 12'hF00;
	mem[12'h321] = 12'hF00;
	mem[12'h322] = 12'hF00;
	mem[12'h323] = 12'hF00;
	mem[12'h324] = 12'hF00;
	mem[12'h325] = 12'hF00;
	mem[12'h326] = 12'hF00;
	mem[12'h327] = 12'hF00;
	mem[12'h328] = 12'hF00;
	mem[12'h329] = 12'hF00;
	mem[12'h32A] = 12'hF00;
	mem[12'h32B] = 12'hF00;
	mem[12'h32C] = 12'hF00;
	mem[12'h32D] = 12'hF00;
	mem[12'h32E] = 12'hF00;
	mem[12'h32F] = 12'hF00;
	mem[12'h330] = 12'hF00;
	mem[12'h331] = 12'hF00;
	mem[12'h332] = 12'hF00;
	mem[12'h333] = 12'hFFF;
	mem[12'h334] = 12'hFFF;
	mem[12'h335] = 12'hFFF;
	mem[12'h336] = 12'hFFF;
	mem[12'h337] = 12'hFFF;
	mem[12'h338] = 12'hFFF;
	mem[12'h339] = 12'hFFF;
	mem[12'h33A] = 12'hFFF;
	mem[12'h33B] = 12'hFFF;
	mem[12'h33C] = 12'hFFF;
	mem[12'h33D] = 12'hFFF;
	mem[12'h33E] = 12'hFFF;
	mem[12'h33F] = 12'hFFF;
	mem[12'h340] = 12'hFFF;
	mem[12'h341] = 12'hFFF;
	mem[12'h342] = 12'hFFF;
	mem[12'h343] = 12'hFFF;
	mem[12'h344] = 12'hFFF;
	mem[12'h345] = 12'hFFF;
	mem[12'h346] = 12'hFFF;
	mem[12'h347] = 12'hFFF;
	mem[12'h348] = 12'hFFF;
	mem[12'h349] = 12'hFFF;
	mem[12'h34A] = 12'hFFF;
	mem[12'h34B] = 12'hFFF;
	mem[12'h34C] = 12'hF00;
	mem[12'h34D] = 12'hF00;
	mem[12'h34E] = 12'hF00;
	mem[12'h34F] = 12'hF00;
	mem[12'h350] = 12'hF00;
	mem[12'h351] = 12'hF00;
	mem[12'h352] = 12'hF00;
	mem[12'h353] = 12'hF00;
	mem[12'h354] = 12'hF00;
	mem[12'h355] = 12'hF00;
	mem[12'h356] = 12'hF00;
	mem[12'h357] = 12'hF00;
	mem[12'h358] = 12'hF00;
	mem[12'h359] = 12'hF00;
	mem[12'h35A] = 12'hF00;
	mem[12'h35B] = 12'hF00;
	mem[12'h35C] = 12'hF00;
	mem[12'h35D] = 12'hF00;
	mem[12'h35E] = 12'hF00;
	mem[12'h35F] = 12'hF00;
	mem[12'h360] = 12'hF00;
	mem[12'h361] = 12'hF00;
	mem[12'h362] = 12'hF00;
	mem[12'h363] = 12'hF00;
	mem[12'h364] = 12'hF00;
	mem[12'h365] = 12'hF00;
	mem[12'h366] = 12'hF00;
	mem[12'h367] = 12'hF00;
	mem[12'h368] = 12'hF00;
	mem[12'h369] = 12'hF00;
	mem[12'h36A] = 12'hF00;
	mem[12'h36B] = 12'hF00;
	mem[12'h36C] = 12'hF00;
	mem[12'h36D] = 12'hF00;
	mem[12'h36E] = 12'hF00;
	mem[12'h36F] = 12'hF00;
	mem[12'h370] = 12'hF00;
	mem[12'h371] = 12'hF00;
	mem[12'h372] = 12'hF00;
	mem[12'h373] = 12'hF00;
	mem[12'h374] = 12'hFFF;
	mem[12'h375] = 12'hFFF;
	mem[12'h376] = 12'hFFF;
	mem[12'h377] = 12'hFFF;
	mem[12'h378] = 12'hFFF;
	mem[12'h379] = 12'hFFF;
	mem[12'h37A] = 12'hFFF;
	mem[12'h37B] = 12'hFFF;
	mem[12'h37C] = 12'hFFF;
	mem[12'h37D] = 12'hFFF;
	mem[12'h37E] = 12'hFFF;
	mem[12'h37F] = 12'hFFF;
	mem[12'h380] = 12'hFFF;
	mem[12'h381] = 12'hFFF;
	mem[12'h382] = 12'hFFF;
	mem[12'h383] = 12'hFFF;
	mem[12'h384] = 12'hFFF;
	mem[12'h385] = 12'hFFF;
	mem[12'h386] = 12'hFFF;
	mem[12'h387] = 12'hFFF;
	mem[12'h388] = 12'hFFF;
	mem[12'h389] = 12'hFFF;
	mem[12'h38A] = 12'hFFF;
	mem[12'h38B] = 12'hF00;
	mem[12'h38C] = 12'hF00;
	mem[12'h38D] = 12'hF00;
	mem[12'h38E] = 12'hF00;
	mem[12'h38F] = 12'hF00;
	mem[12'h390] = 12'hF00;
	mem[12'h391] = 12'hF00;
	mem[12'h392] = 12'hF00;
	mem[12'h393] = 12'hF00;
	mem[12'h394] = 12'hF00;
	mem[12'h395] = 12'hF00;
	mem[12'h396] = 12'hF00;
	mem[12'h397] = 12'hF00;
	mem[12'h398] = 12'hF00;
	mem[12'h399] = 12'hF00;
	mem[12'h39A] = 12'hF00;
	mem[12'h39B] = 12'hF00;
	mem[12'h39C] = 12'hF00;
	mem[12'h39D] = 12'hF00;
	mem[12'h39E] = 12'hF00;
	mem[12'h39F] = 12'hF00;
	mem[12'h3A0] = 12'hF00;
	mem[12'h3A1] = 12'hF00;
	mem[12'h3A2] = 12'hF00;
	mem[12'h3A3] = 12'hF00;
	mem[12'h3A4] = 12'hF00;
	mem[12'h3A5] = 12'hF00;
	mem[12'h3A6] = 12'hF00;
	mem[12'h3A7] = 12'hF00;
	mem[12'h3A8] = 12'hF00;
	mem[12'h3A9] = 12'hF00;
	mem[12'h3AA] = 12'hF00;
	mem[12'h3AB] = 12'hF00;
	mem[12'h3AC] = 12'hF00;
	mem[12'h3AD] = 12'hF00;
	mem[12'h3AE] = 12'hF00;
	mem[12'h3AF] = 12'hF00;
	mem[12'h3B0] = 12'hF00;
	mem[12'h3B1] = 12'hF00;
	mem[12'h3B2] = 12'hF00;
	mem[12'h3B3] = 12'hF00;
	mem[12'h3B4] = 12'hF00;
	mem[12'h3B5] = 12'hFFF;
	mem[12'h3B6] = 12'hFFF;
	mem[12'h3B7] = 12'hFFF;
	mem[12'h3B8] = 12'hFFF;
	mem[12'h3B9] = 12'hFFF;
	mem[12'h3BA] = 12'hFFF;
	mem[12'h3BB] = 12'hFFF;
	mem[12'h3BC] = 12'hFFF;
	mem[12'h3BD] = 12'hFFF;
	mem[12'h3BE] = 12'hFFF;
	mem[12'h3BF] = 12'hFFF;
	mem[12'h3C0] = 12'hFFF;
	mem[12'h3C1] = 12'hFFF;
	mem[12'h3C2] = 12'hFFF;
	mem[12'h3C3] = 12'hFFF;
	mem[12'h3C4] = 12'hFFF;
	mem[12'h3C5] = 12'hFFF;
	mem[12'h3C6] = 12'hFFF;
	mem[12'h3C7] = 12'hFFF;
	mem[12'h3C8] = 12'hFFF;
	mem[12'h3C9] = 12'hFFF;
	mem[12'h3CA] = 12'hFFF;
	mem[12'h3CB] = 12'hE22;
	mem[12'h3CC] = 12'hF00;
	mem[12'h3CD] = 12'hF00;
	mem[12'h3CE] = 12'hF00;
	mem[12'h3CF] = 12'hF00;
	mem[12'h3D0] = 12'hF00;
	mem[12'h3D1] = 12'hF00;
	mem[12'h3D2] = 12'hF00;
	mem[12'h3D3] = 12'hF00;
	mem[12'h3D4] = 12'hF00;
	mem[12'h3D5] = 12'hF00;
	mem[12'h3D6] = 12'hF00;
	mem[12'h3D7] = 12'hF00;
	mem[12'h3D8] = 12'hF00;
	mem[12'h3D9] = 12'hF00;
	mem[12'h3DA] = 12'hF00;
	mem[12'h3DB] = 12'hF00;
	mem[12'h3DC] = 12'hF00;
	mem[12'h3DD] = 12'hF00;
	mem[12'h3DE] = 12'hF00;
	mem[12'h3DF] = 12'hF00;
	mem[12'h3E0] = 12'hF00;
	mem[12'h3E1] = 12'hF00;
	mem[12'h3E2] = 12'hF00;
	mem[12'h3E3] = 12'hF00;
	mem[12'h3E4] = 12'hF00;
	mem[12'h3E5] = 12'hF00;
	mem[12'h3E6] = 12'hF00;
	mem[12'h3E7] = 12'hF00;
	mem[12'h3E8] = 12'hF00;
	mem[12'h3E9] = 12'hF00;
	mem[12'h3EA] = 12'hF00;
	mem[12'h3EB] = 12'hF00;
	mem[12'h3EC] = 12'hF00;
	mem[12'h3ED] = 12'hF00;
	mem[12'h3EE] = 12'hF00;
	mem[12'h3EF] = 12'hF00;
	mem[12'h3F0] = 12'hF00;
	mem[12'h3F1] = 12'hF00;
	mem[12'h3F2] = 12'hF00;
	mem[12'h3F3] = 12'hF00;
	mem[12'h3F4] = 12'hE22;
	mem[12'h3F5] = 12'hFFF;
	mem[12'h3F6] = 12'hFFF;
	mem[12'h3F7] = 12'hFFF;
	mem[12'h3F8] = 12'hFFF;
	mem[12'h3F9] = 12'hFFF;
	mem[12'h3FA] = 12'hFFF;
	mem[12'h3FB] = 12'hFFF;
	mem[12'h3FC] = 12'hFFF;
	mem[12'h3FD] = 12'hFFF;
	mem[12'h3FE] = 12'hFFF;
	mem[12'h3FF] = 12'hFFF;
	mem[12'h400] = 12'hFFF;
	mem[12'h401] = 12'hFFF;
	mem[12'h402] = 12'hFFF;
	mem[12'h403] = 12'hFFF;
	mem[12'h404] = 12'hFFF;
	mem[12'h405] = 12'hFFF;
	mem[12'h406] = 12'hFFF;
	mem[12'h407] = 12'hFFF;
	mem[12'h408] = 12'hFFF;
	mem[12'h409] = 12'hFFF;
	mem[12'h40A] = 12'hF00;
	mem[12'h40B] = 12'hF00;
	mem[12'h40C] = 12'hF00;
	mem[12'h40D] = 12'hF00;
	mem[12'h40E] = 12'hF00;
	mem[12'h40F] = 12'hF00;
	mem[12'h410] = 12'hF00;
	mem[12'h411] = 12'hF00;
	mem[12'h412] = 12'hF00;
	mem[12'h413] = 12'hF00;
	mem[12'h414] = 12'hF00;
	mem[12'h415] = 12'hF00;
	mem[12'h416] = 12'hF00;
	mem[12'h417] = 12'hF00;
	mem[12'h418] = 12'hF00;
	mem[12'h419] = 12'hF00;
	mem[12'h41A] = 12'hF00;
	mem[12'h41B] = 12'hF00;
	mem[12'h41C] = 12'hF00;
	mem[12'h41D] = 12'hF00;
	mem[12'h41E] = 12'hF00;
	mem[12'h41F] = 12'hF00;
	mem[12'h420] = 12'hF00;
	mem[12'h421] = 12'hF00;
	mem[12'h422] = 12'hF00;
	mem[12'h423] = 12'hF00;
	mem[12'h424] = 12'hF00;
	mem[12'h425] = 12'hF00;
	mem[12'h426] = 12'hF00;
	mem[12'h427] = 12'hF00;
	mem[12'h428] = 12'hF00;
	mem[12'h429] = 12'hF00;
	mem[12'h42A] = 12'hF00;
	mem[12'h42B] = 12'hF00;
	mem[12'h42C] = 12'hF00;
	mem[12'h42D] = 12'hF00;
	mem[12'h42E] = 12'hF00;
	mem[12'h42F] = 12'hF00;
	mem[12'h430] = 12'hF00;
	mem[12'h431] = 12'hF00;
	mem[12'h432] = 12'hF00;
	mem[12'h433] = 12'hF00;
	mem[12'h434] = 12'hF00;
	mem[12'h435] = 12'hE22;
	mem[12'h436] = 12'hFFF;
	mem[12'h437] = 12'hFFF;
	mem[12'h438] = 12'hFFF;
	mem[12'h439] = 12'hFFF;
	mem[12'h43A] = 12'hFFF;
	mem[12'h43B] = 12'hFFF;
	mem[12'h43C] = 12'hFFF;
	mem[12'h43D] = 12'hFFF;
	mem[12'h43E] = 12'hFFF;
	mem[12'h43F] = 12'hFFF;
	mem[12'h440] = 12'hFFF;
	mem[12'h441] = 12'hFFF;
	mem[12'h442] = 12'hFFF;
	mem[12'h443] = 12'hFFF;
	mem[12'h444] = 12'hFFF;
	mem[12'h445] = 12'hFFF;
	mem[12'h446] = 12'hFFF;
	mem[12'h447] = 12'hFFF;
	mem[12'h448] = 12'hFFF;
	mem[12'h449] = 12'hFFF;
	mem[12'h44A] = 12'hF00;
	mem[12'h44B] = 12'hF00;
	mem[12'h44C] = 12'hF00;
	mem[12'h44D] = 12'hF00;
	mem[12'h44E] = 12'hF00;
	mem[12'h44F] = 12'hF00;
	mem[12'h450] = 12'hF00;
	mem[12'h451] = 12'hF00;
	mem[12'h452] = 12'hF00;
	mem[12'h453] = 12'hF00;
	mem[12'h454] = 12'hF00;
	mem[12'h455] = 12'hF00;
	mem[12'h456] = 12'hF00;
	mem[12'h457] = 12'hF00;
	mem[12'h458] = 12'hF00;
	mem[12'h459] = 12'hF00;
	mem[12'h45A] = 12'hF00;
	mem[12'h45B] = 12'hF00;
	mem[12'h45C] = 12'hF00;
	mem[12'h45D] = 12'hF00;
	mem[12'h45E] = 12'hF00;
	mem[12'h45F] = 12'hF00;
	mem[12'h460] = 12'hF00;
	mem[12'h461] = 12'hF00;
	mem[12'h462] = 12'hF00;
	mem[12'h463] = 12'hF00;
	mem[12'h464] = 12'hF00;
	mem[12'h465] = 12'hF00;
	mem[12'h466] = 12'hF00;
	mem[12'h467] = 12'hF00;
	mem[12'h468] = 12'hF00;
	mem[12'h469] = 12'hF00;
	mem[12'h46A] = 12'hF00;
	mem[12'h46B] = 12'hF00;
	mem[12'h46C] = 12'hF00;
	mem[12'h46D] = 12'hF00;
	mem[12'h46E] = 12'hF00;
	mem[12'h46F] = 12'hF00;
	mem[12'h470] = 12'hF00;
	mem[12'h471] = 12'hF00;
	mem[12'h472] = 12'hF00;
	mem[12'h473] = 12'hF00;
	mem[12'h474] = 12'hF00;
	mem[12'h475] = 12'hF00;
	mem[12'h476] = 12'hFFF;
	mem[12'h477] = 12'hFFF;
	mem[12'h478] = 12'hFFF;
	mem[12'h479] = 12'hFFF;
	mem[12'h47A] = 12'hFFF;
	mem[12'h47B] = 12'hFFF;
	mem[12'h47C] = 12'hFFF;
	mem[12'h47D] = 12'hFFF;
	mem[12'h47E] = 12'hFFF;
	mem[12'h47F] = 12'hFFF;
	mem[12'h480] = 12'hFFF;
	mem[12'h481] = 12'hFFF;
	mem[12'h482] = 12'hFFF;
	mem[12'h483] = 12'hFFF;
	mem[12'h484] = 12'hFFF;
	mem[12'h485] = 12'hFFF;
	mem[12'h486] = 12'hFFF;
	mem[12'h487] = 12'hFFF;
	mem[12'h488] = 12'hFFF;
	mem[12'h489] = 12'hE22;
	mem[12'h48A] = 12'hF00;
	mem[12'h48B] = 12'hF00;
	mem[12'h48C] = 12'hF00;
	mem[12'h48D] = 12'hF00;
	mem[12'h48E] = 12'hF00;
	mem[12'h48F] = 12'hF00;
	mem[12'h490] = 12'hF00;
	mem[12'h491] = 12'hF00;
	mem[12'h492] = 12'hF00;
	mem[12'h493] = 12'hF00;
	mem[12'h494] = 12'hF00;
	mem[12'h495] = 12'hF00;
	mem[12'h496] = 12'hF00;
	mem[12'h497] = 12'hF00;
	mem[12'h498] = 12'hF00;
	mem[12'h499] = 12'hF00;
	mem[12'h49A] = 12'hF00;
	mem[12'h49B] = 12'hF00;
	mem[12'h49C] = 12'hF00;
	mem[12'h49D] = 12'hF00;
	mem[12'h49E] = 12'hF00;
	mem[12'h49F] = 12'hF00;
	mem[12'h4A0] = 12'hF00;
	mem[12'h4A1] = 12'hF00;
	mem[12'h4A2] = 12'hF00;
	mem[12'h4A3] = 12'hF00;
	mem[12'h4A4] = 12'hF00;
	mem[12'h4A5] = 12'hF00;
	mem[12'h4A6] = 12'hF00;
	mem[12'h4A7] = 12'hF00;
	mem[12'h4A8] = 12'hF00;
	mem[12'h4A9] = 12'hF00;
	mem[12'h4AA] = 12'hF00;
	mem[12'h4AB] = 12'hF00;
	mem[12'h4AC] = 12'hF00;
	mem[12'h4AD] = 12'hF00;
	mem[12'h4AE] = 12'hF00;
	mem[12'h4AF] = 12'hF00;
	mem[12'h4B0] = 12'hF00;
	mem[12'h4B1] = 12'hF00;
	mem[12'h4B2] = 12'hF00;
	mem[12'h4B3] = 12'hF00;
	mem[12'h4B4] = 12'hF00;
	mem[12'h4B5] = 12'hF00;
	mem[12'h4B6] = 12'hE22;
	mem[12'h4B7] = 12'hFFF;
	mem[12'h4B8] = 12'hFFF;
	mem[12'h4B9] = 12'hFFF;
	mem[12'h4BA] = 12'hFFF;
	mem[12'h4BB] = 12'hFFF;
	mem[12'h4BC] = 12'hFFF;
	mem[12'h4BD] = 12'hFFF;
	mem[12'h4BE] = 12'hFFF;
	mem[12'h4BF] = 12'hFFF;
	mem[12'h4C0] = 12'hFFF;
	mem[12'h4C1] = 12'hFFF;
	mem[12'h4C2] = 12'hFFF;
	mem[12'h4C3] = 12'hFFF;
	mem[12'h4C4] = 12'hFFF;
	mem[12'h4C5] = 12'hFFF;
	mem[12'h4C6] = 12'hFFF;
	mem[12'h4C7] = 12'hFFF;
	mem[12'h4C8] = 12'hFFF;
	mem[12'h4C9] = 12'hF00;
	mem[12'h4CA] = 12'hF00;
	mem[12'h4CB] = 12'hF00;
	mem[12'h4CC] = 12'hF00;
	mem[12'h4CD] = 12'hF00;
	mem[12'h4CE] = 12'hF00;
	mem[12'h4CF] = 12'hF00;
	mem[12'h4D0] = 12'hF00;
	mem[12'h4D1] = 12'hF00;
	mem[12'h4D2] = 12'hF00;
	mem[12'h4D3] = 12'hF00;
	mem[12'h4D4] = 12'hF00;
	mem[12'h4D5] = 12'hF00;
	mem[12'h4D6] = 12'hF00;
	mem[12'h4D7] = 12'hF00;
	mem[12'h4D8] = 12'hF00;
	mem[12'h4D9] = 12'hF00;
	mem[12'h4DA] = 12'hF00;
	mem[12'h4DB] = 12'hF00;
	mem[12'h4DC] = 12'hF00;
	mem[12'h4DD] = 12'hF00;
	mem[12'h4DE] = 12'hF00;
	mem[12'h4DF] = 12'hF00;
	mem[12'h4E0] = 12'hF00;
	mem[12'h4E1] = 12'hF00;
	mem[12'h4E2] = 12'hF00;
	mem[12'h4E3] = 12'hF00;
	mem[12'h4E4] = 12'hF00;
	mem[12'h4E5] = 12'hF00;
	mem[12'h4E6] = 12'hF00;
	mem[12'h4E7] = 12'hF00;
	mem[12'h4E8] = 12'hF00;
	mem[12'h4E9] = 12'hF00;
	mem[12'h4EA] = 12'hF00;
	mem[12'h4EB] = 12'hF00;
	mem[12'h4EC] = 12'hF00;
	mem[12'h4ED] = 12'hF00;
	mem[12'h4EE] = 12'hF00;
	mem[12'h4EF] = 12'hF00;
	mem[12'h4F0] = 12'hF00;
	mem[12'h4F1] = 12'hF00;
	mem[12'h4F2] = 12'hF00;
	mem[12'h4F3] = 12'hF00;
	mem[12'h4F4] = 12'hF00;
	mem[12'h4F5] = 12'hF00;
	mem[12'h4F6] = 12'hF00;
	mem[12'h4F7] = 12'hFFF;
	mem[12'h4F8] = 12'hFFF;
	mem[12'h4F9] = 12'hFFF;
	mem[12'h4FA] = 12'hFFF;
	mem[12'h4FB] = 12'hFFF;
	mem[12'h4FC] = 12'hFFF;
	mem[12'h4FD] = 12'hFFF;
	mem[12'h4FE] = 12'hFFF;
	mem[12'h4FF] = 12'hFFF;
	mem[12'h500] = 12'hFFF;
	mem[12'h501] = 12'hFFF;
	mem[12'h502] = 12'hFFF;
	mem[12'h503] = 12'hFFF;
	mem[12'h504] = 12'hFFF;
	mem[12'h505] = 12'hFFF;
	mem[12'h506] = 12'hFFF;
	mem[12'h507] = 12'hFFF;
	mem[12'h508] = 12'hF00;
	mem[12'h509] = 12'hF00;
	mem[12'h50A] = 12'hF00;
	mem[12'h50B] = 12'hF00;
	mem[12'h50C] = 12'hF00;
	mem[12'h50D] = 12'hF00;
	mem[12'h50E] = 12'hF00;
	mem[12'h50F] = 12'hF00;
	mem[12'h510] = 12'hF00;
	mem[12'h511] = 12'hF00;
	mem[12'h512] = 12'hF00;
	mem[12'h513] = 12'hF00;
	mem[12'h514] = 12'hF00;
	mem[12'h515] = 12'hF00;
	mem[12'h516] = 12'hF00;
	mem[12'h517] = 12'hE22;
	mem[12'h518] = 12'hF00;
	mem[12'h519] = 12'hFFF;
	mem[12'h51A] = 12'hFFF;
	mem[12'h51B] = 12'hFFF;
	mem[12'h51C] = 12'hF00;
	mem[12'h51D] = 12'hE22;
	mem[12'h51E] = 12'hF00;
	mem[12'h51F] = 12'hF00;
	mem[12'h520] = 12'hF00;
	mem[12'h521] = 12'hF00;
	mem[12'h522] = 12'hF00;
	mem[12'h523] = 12'hF00;
	mem[12'h524] = 12'hF00;
	mem[12'h525] = 12'hF00;
	mem[12'h526] = 12'hF00;
	mem[12'h527] = 12'hF00;
	mem[12'h528] = 12'hF00;
	mem[12'h529] = 12'hF00;
	mem[12'h52A] = 12'hF00;
	mem[12'h52B] = 12'hF00;
	mem[12'h52C] = 12'hE22;
	mem[12'h52D] = 12'hF00;
	mem[12'h52E] = 12'hFFF;
	mem[12'h52F] = 12'hFFF;
	mem[12'h530] = 12'hF00;
	mem[12'h531] = 12'hF00;
	mem[12'h532] = 12'hF00;
	mem[12'h533] = 12'hF00;
	mem[12'h534] = 12'hF00;
	mem[12'h535] = 12'hF00;
	mem[12'h536] = 12'hF00;
	mem[12'h537] = 12'hF00;
	mem[12'h538] = 12'hFFF;
	mem[12'h539] = 12'hFFF;
	mem[12'h53A] = 12'hFFF;
	mem[12'h53B] = 12'hFFF;
	mem[12'h53C] = 12'hFFF;
	mem[12'h53D] = 12'hFFF;
	mem[12'h53E] = 12'hFFF;
	mem[12'h53F] = 12'hFFF;
	mem[12'h540] = 12'hFFF;
	mem[12'h541] = 12'hFFF;
	mem[12'h542] = 12'hFFF;
	mem[12'h543] = 12'hFFF;
	mem[12'h544] = 12'hFFF;
	mem[12'h545] = 12'hFFF;
	mem[12'h546] = 12'hFFF;
	mem[12'h547] = 12'hFFF;
	mem[12'h548] = 12'hE22;
	mem[12'h549] = 12'hF00;
	mem[12'h54A] = 12'hF00;
	mem[12'h54B] = 12'hF00;
	mem[12'h54C] = 12'hF00;
	mem[12'h54D] = 12'hF00;
	mem[12'h54E] = 12'hF00;
	mem[12'h54F] = 12'hF00;
	mem[12'h550] = 12'hF00;
	mem[12'h551] = 12'hF00;
	mem[12'h552] = 12'hF00;
	mem[12'h553] = 12'hF00;
	mem[12'h554] = 12'hF00;
	mem[12'h555] = 12'hF00;
	mem[12'h556] = 12'hE22;
	mem[12'h557] = 12'hFFF;
	mem[12'h558] = 12'hFFF;
	mem[12'h559] = 12'hFFF;
	mem[12'h55A] = 12'hFFF;
	mem[12'h55B] = 12'hFFF;
	mem[12'h55C] = 12'hFFF;
	mem[12'h55D] = 12'hFFF;
	mem[12'h55E] = 12'hF00;
	mem[12'h55F] = 12'hF00;
	mem[12'h560] = 12'hF00;
	mem[12'h561] = 12'hF00;
	mem[12'h562] = 12'hF00;
	mem[12'h563] = 12'hF00;
	mem[12'h564] = 12'hF00;
	mem[12'h565] = 12'hF00;
	mem[12'h566] = 12'hF00;
	mem[12'h567] = 12'hF00;
	mem[12'h568] = 12'hF00;
	mem[12'h569] = 12'hF00;
	mem[12'h56A] = 12'hE22;
	mem[12'h56B] = 12'hFFF;
	mem[12'h56C] = 12'hFFF;
	mem[12'h56D] = 12'hFFF;
	mem[12'h56E] = 12'hFFF;
	mem[12'h56F] = 12'hFFF;
	mem[12'h570] = 12'hFFF;
	mem[12'h571] = 12'hFFF;
	mem[12'h572] = 12'hFFF;
	mem[12'h573] = 12'hE22;
	mem[12'h574] = 12'hF00;
	mem[12'h575] = 12'hF00;
	mem[12'h576] = 12'hF00;
	mem[12'h577] = 12'hE22;
	mem[12'h578] = 12'hFFF;
	mem[12'h579] = 12'hFFF;
	mem[12'h57A] = 12'hFFF;
	mem[12'h57B] = 12'hFFF;
	mem[12'h57C] = 12'hFFF;
	mem[12'h57D] = 12'hFFF;
	mem[12'h57E] = 12'hFFF;
	mem[12'h57F] = 12'hFFF;
	mem[12'h580] = 12'hFFF;
	mem[12'h581] = 12'hFFF;
	mem[12'h582] = 12'hFFF;
	mem[12'h583] = 12'hFFF;
	mem[12'h584] = 12'hFFF;
	mem[12'h585] = 12'hFFF;
	mem[12'h586] = 12'hFFF;
	mem[12'h587] = 12'hFFF;
	mem[12'h588] = 12'hF00;
	mem[12'h589] = 12'hF00;
	mem[12'h58A] = 12'hF00;
	mem[12'h58B] = 12'hF00;
	mem[12'h58C] = 12'hF00;
	mem[12'h58D] = 12'hF00;
	mem[12'h58E] = 12'hF00;
	mem[12'h58F] = 12'hF00;
	mem[12'h590] = 12'hF00;
	mem[12'h591] = 12'hF00;
	mem[12'h592] = 12'hF00;
	mem[12'h593] = 12'hF00;
	mem[12'h594] = 12'hF00;
	mem[12'h595] = 12'hF00;
	mem[12'h596] = 12'hFFF;
	mem[12'h597] = 12'hFFF;
	mem[12'h598] = 12'hFFF;
	mem[12'h599] = 12'hFFF;
	mem[12'h59A] = 12'hFFF;
	mem[12'h59B] = 12'hFFF;
	mem[12'h59C] = 12'hFFF;
	mem[12'h59D] = 12'hFFF;
	mem[12'h59E] = 12'hFFF;
	mem[12'h59F] = 12'hF00;
	mem[12'h5A0] = 12'hF00;
	mem[12'h5A1] = 12'hF00;
	mem[12'h5A2] = 12'hF00;
	mem[12'h5A3] = 12'hF00;
	mem[12'h5A4] = 12'hF00;
	mem[12'h5A5] = 12'hF00;
	mem[12'h5A6] = 12'hF00;
	mem[12'h5A7] = 12'hF00;
	mem[12'h5A8] = 12'hF00;
	mem[12'h5A9] = 12'hE22;
	mem[12'h5AA] = 12'hFFF;
	mem[12'h5AB] = 12'hFFF;
	mem[12'h5AC] = 12'hFFF;
	mem[12'h5AD] = 12'hFFF;
	mem[12'h5AE] = 12'hFFF;
	mem[12'h5AF] = 12'hFFF;
	mem[12'h5B0] = 12'hFFF;
	mem[12'h5B1] = 12'hFFF;
	mem[12'h5B2] = 12'hFFF;
	mem[12'h5B3] = 12'hFFF;
	mem[12'h5B4] = 12'hE22;
	mem[12'h5B5] = 12'hF00;
	mem[12'h5B6] = 12'hF00;
	mem[12'h5B7] = 12'hF00;
	mem[12'h5B8] = 12'hFFF;
	mem[12'h5B9] = 12'hFFF;
	mem[12'h5BA] = 12'hFFF;
	mem[12'h5BB] = 12'hFFF;
	mem[12'h5BC] = 12'hFFF;
	mem[12'h5BD] = 12'hFFF;
	mem[12'h5BE] = 12'hFFF;
	mem[12'h5BF] = 12'hFFF;
	mem[12'h5C0] = 12'hFFF;
	mem[12'h5C1] = 12'hFFF;
	mem[12'h5C2] = 12'hFFF;
	mem[12'h5C3] = 12'hFFF;
	mem[12'h5C4] = 12'hFFF;
	mem[12'h5C5] = 12'hFFF;
	mem[12'h5C6] = 12'hFFF;
	mem[12'h5C7] = 12'hFFF;
	mem[12'h5C8] = 12'hF00;
	mem[12'h5C9] = 12'hF00;
	mem[12'h5CA] = 12'hF00;
	mem[12'h5CB] = 12'hF00;
	mem[12'h5CC] = 12'hF00;
	mem[12'h5CD] = 12'hF00;
	mem[12'h5CE] = 12'hF00;
	mem[12'h5CF] = 12'hF00;
	mem[12'h5D0] = 12'hF00;
	mem[12'h5D1] = 12'hF00;
	mem[12'h5D2] = 12'hF00;
	mem[12'h5D3] = 12'hF00;
	mem[12'h5D4] = 12'hE22;
	mem[12'h5D5] = 12'hFFF;
	mem[12'h5D6] = 12'hFFF;
	mem[12'h5D7] = 12'hFFF;
	mem[12'h5D8] = 12'hFFF;
	mem[12'h5D9] = 12'hFFF;
	mem[12'h5DA] = 12'hFFF;
	mem[12'h5DB] = 12'hFFF;
	mem[12'h5DC] = 12'hFFF;
	mem[12'h5DD] = 12'hFFF;
	mem[12'h5DE] = 12'hFFF;
	mem[12'h5DF] = 12'hFFF;
	mem[12'h5E0] = 12'hF00;
	mem[12'h5E1] = 12'hF00;
	mem[12'h5E2] = 12'hF00;
	mem[12'h5E3] = 12'hF00;
	mem[12'h5E4] = 12'hF00;
	mem[12'h5E5] = 12'hF00;
	mem[12'h5E6] = 12'hF00;
	mem[12'h5E7] = 12'hF00;
	mem[12'h5E8] = 12'hF00;
	mem[12'h5E9] = 12'hFFF;
	mem[12'h5EA] = 12'hFFF;
	mem[12'h5EB] = 12'hFFF;
	mem[12'h5EC] = 12'hFFF;
	mem[12'h5ED] = 12'hFFF;
	mem[12'h5EE] = 12'hFFF;
	mem[12'h5EF] = 12'hFFF;
	mem[12'h5F0] = 12'hFFF;
	mem[12'h5F1] = 12'hFFF;
	mem[12'h5F2] = 12'hFFF;
	mem[12'h5F3] = 12'hFFF;
	mem[12'h5F4] = 12'hFFF;
	mem[12'h5F5] = 12'hF00;
	mem[12'h5F6] = 12'hF00;
	mem[12'h5F7] = 12'hF00;
	mem[12'h5F8] = 12'hFFF;
	mem[12'h5F9] = 12'hFFF;
	mem[12'h5FA] = 12'hFFF;
	mem[12'h5FB] = 12'hFFF;
	mem[12'h5FC] = 12'hFFF;
	mem[12'h5FD] = 12'hFFF;
	mem[12'h5FE] = 12'hFFF;
	mem[12'h5FF] = 12'hFFF;
	mem[12'h600] = 12'hFFF;
	mem[12'h601] = 12'hFFF;
	mem[12'h602] = 12'hFFF;
	mem[12'h603] = 12'hFFF;
	mem[12'h604] = 12'hFFF;
	mem[12'h605] = 12'hFFF;
	mem[12'h606] = 12'hFFF;
	mem[12'h607] = 12'hF00;
	mem[12'h608] = 12'hF00;
	mem[12'h609] = 12'hF00;
	mem[12'h60A] = 12'hF00;
	mem[12'h60B] = 12'hF00;
	mem[12'h60C] = 12'hF00;
	mem[12'h60D] = 12'hF00;
	mem[12'h60E] = 12'hF00;
	mem[12'h60F] = 12'hF00;
	mem[12'h610] = 12'hF00;
	mem[12'h611] = 12'hF00;
	mem[12'h612] = 12'hF00;
	mem[12'h613] = 12'hF00;
	mem[12'h614] = 12'hF00;
	mem[12'h615] = 12'hFFF;
	mem[12'h616] = 12'hFFF;
	mem[12'h617] = 12'hFFF;
	mem[12'h618] = 12'hFFF;
	mem[12'h619] = 12'hFFF;
	mem[12'h61A] = 12'hFFF;
	mem[12'h61B] = 12'h01C;
	mem[12'h61C] = 12'h01C;
	mem[12'h61D] = 12'h01C;
	mem[12'h61E] = 12'h01C;
	mem[12'h61F] = 12'h01C;
	mem[12'h620] = 12'hFFF;
	mem[12'h621] = 12'hF00;
	mem[12'h622] = 12'hF00;
	mem[12'h623] = 12'hF00;
	mem[12'h624] = 12'hF00;
	mem[12'h625] = 12'hF00;
	mem[12'h626] = 12'hF00;
	mem[12'h627] = 12'hF00;
	mem[12'h628] = 12'hE22;
	mem[12'h629] = 12'hFFF;
	mem[12'h62A] = 12'hFFF;
	mem[12'h62B] = 12'hFFF;
	mem[12'h62C] = 12'hFFF;
	mem[12'h62D] = 12'hFFF;
	mem[12'h62E] = 12'hFFF;
	mem[12'h62F] = 12'h01C;
	mem[12'h630] = 12'h01C;
	mem[12'h631] = 12'h01C;
	mem[12'h632] = 12'h01C;
	mem[12'h633] = 12'h01C;
	mem[12'h634] = 12'hFFF;
	mem[12'h635] = 12'hF00;
	mem[12'h636] = 12'hF00;
	mem[12'h637] = 12'hF00;
	mem[12'h638] = 12'hF00;
	mem[12'h639] = 12'hFFF;
	mem[12'h63A] = 12'hFFF;
	mem[12'h63B] = 12'hFFF;
	mem[12'h63C] = 12'hFFF;
	mem[12'h63D] = 12'hFFF;
	mem[12'h63E] = 12'hFFF;
	mem[12'h63F] = 12'hFFF;
	mem[12'h640] = 12'hFFF;
	mem[12'h641] = 12'hFFF;
	mem[12'h642] = 12'hFFF;
	mem[12'h643] = 12'hFFF;
	mem[12'h644] = 12'hFFF;
	mem[12'h645] = 12'hFFF;
	mem[12'h646] = 12'hFFF;
	mem[12'h647] = 12'hF00;
	mem[12'h648] = 12'hF00;
	mem[12'h649] = 12'hF00;
	mem[12'h64A] = 12'hF00;
	mem[12'h64B] = 12'hF00;
	mem[12'h64C] = 12'hF00;
	mem[12'h64D] = 12'hF00;
	mem[12'h64E] = 12'hF00;
	mem[12'h64F] = 12'hF00;
	mem[12'h650] = 12'hF00;
	mem[12'h651] = 12'hF00;
	mem[12'h652] = 12'hF00;
	mem[12'h653] = 12'hF00;
	mem[12'h654] = 12'hFFF;
	mem[12'h655] = 12'hFFF;
	mem[12'h656] = 12'hFFF;
	mem[12'h657] = 12'hFFF;
	mem[12'h658] = 12'hFFF;
	mem[12'h659] = 12'hFFF;
	mem[12'h65A] = 12'h01C;
	mem[12'h65B] = 12'h01C;
	mem[12'h65C] = 12'h00C;
	mem[12'h65D] = 12'h00C;
	mem[12'h65E] = 12'h00C;
	mem[12'h65F] = 12'h01C;
	mem[12'h660] = 12'hFFF;
	mem[12'h661] = 12'hE22;
	mem[12'h662] = 12'hF00;
	mem[12'h663] = 12'hF00;
	mem[12'h664] = 12'hF00;
	mem[12'h665] = 12'hF00;
	mem[12'h666] = 12'hF00;
	mem[12'h667] = 12'hF00;
	mem[12'h668] = 12'hF00;
	mem[12'h669] = 12'hFFF;
	mem[12'h66A] = 12'hFFF;
	mem[12'h66B] = 12'hFFF;
	mem[12'h66C] = 12'hFFF;
	mem[12'h66D] = 12'hFFF;
	mem[12'h66E] = 12'hFFF;
	mem[12'h66F] = 12'h01C;
	mem[12'h670] = 12'h00C;
	mem[12'h671] = 12'h00C;
	mem[12'h672] = 12'h00C;
	mem[12'h673] = 12'h01C;
	mem[12'h674] = 12'h01C;
	mem[12'h675] = 12'hF00;
	mem[12'h676] = 12'hF00;
	mem[12'h677] = 12'hF00;
	mem[12'h678] = 12'hF00;
	mem[12'h679] = 12'hFFF;
	mem[12'h67A] = 12'hFFF;
	mem[12'h67B] = 12'hFFF;
	mem[12'h67C] = 12'hFFF;
	mem[12'h67D] = 12'hFFF;
	mem[12'h67E] = 12'hFFF;
	mem[12'h67F] = 12'hFFF;
	mem[12'h680] = 12'hFFF;
	mem[12'h681] = 12'hFFF;
	mem[12'h682] = 12'hFFF;
	mem[12'h683] = 12'hFFF;
	mem[12'h684] = 12'hFFF;
	mem[12'h685] = 12'hFFF;
	mem[12'h686] = 12'hFFF;
	mem[12'h687] = 12'hF00;
	mem[12'h688] = 12'hF00;
	mem[12'h689] = 12'hF00;
	mem[12'h68A] = 12'hF00;
	mem[12'h68B] = 12'hF00;
	mem[12'h68C] = 12'hF00;
	mem[12'h68D] = 12'hF00;
	mem[12'h68E] = 12'hF00;
	mem[12'h68F] = 12'hF00;
	mem[12'h690] = 12'hF00;
	mem[12'h691] = 12'hF00;
	mem[12'h692] = 12'hF00;
	mem[12'h693] = 12'hF00;
	mem[12'h694] = 12'hFFF;
	mem[12'h695] = 12'hFFF;
	mem[12'h696] = 12'hFFF;
	mem[12'h697] = 12'hFFF;
	mem[12'h698] = 12'hFFF;
	mem[12'h699] = 12'hFFF;
	mem[12'h69A] = 12'h01C;
	mem[12'h69B] = 12'h00C;
	mem[12'h69C] = 12'h00C;
	mem[12'h69D] = 12'h00C;
	mem[12'h69E] = 12'h00C;
	mem[12'h69F] = 12'h01C;
	mem[12'h6A0] = 12'h01C;
	mem[12'h6A1] = 12'hE22;
	mem[12'h6A2] = 12'hF00;
	mem[12'h6A3] = 12'hF00;
	mem[12'h6A4] = 12'hF00;
	mem[12'h6A5] = 12'hF00;
	mem[12'h6A6] = 12'hF00;
	mem[12'h6A7] = 12'hF00;
	mem[12'h6A8] = 12'hFFF;
	mem[12'h6A9] = 12'hFFF;
	mem[12'h6AA] = 12'hFFF;
	mem[12'h6AB] = 12'hFFF;
	mem[12'h6AC] = 12'hFFF;
	mem[12'h6AD] = 12'hFFF;
	mem[12'h6AE] = 12'h01C;
	mem[12'h6AF] = 12'h01C;
	mem[12'h6B0] = 12'h00C;
	mem[12'h6B1] = 12'h00C;
	mem[12'h6B2] = 12'h00C;
	mem[12'h6B3] = 12'h00C;
	mem[12'h6B4] = 12'h01C;
	mem[12'h6B5] = 12'hFFF;
	mem[12'h6B6] = 12'hF00;
	mem[12'h6B7] = 12'hF00;
	mem[12'h6B8] = 12'hF00;
	mem[12'h6B9] = 12'hFFF;
	mem[12'h6BA] = 12'hFFF;
	mem[12'h6BB] = 12'hFFF;
	mem[12'h6BC] = 12'hFFF;
	mem[12'h6BD] = 12'hFFF;
	mem[12'h6BE] = 12'hFFF;
	mem[12'h6BF] = 12'hFFF;
	mem[12'h6C0] = 12'hFFF;
	mem[12'h6C1] = 12'hFFF;
	mem[12'h6C2] = 12'hFFF;
	mem[12'h6C3] = 12'hFFF;
	mem[12'h6C4] = 12'hFFF;
	mem[12'h6C5] = 12'hFFF;
	mem[12'h6C6] = 12'hFFF;
	mem[12'h6C7] = 12'hE22;
	mem[12'h6C8] = 12'hF00;
	mem[12'h6C9] = 12'hF00;
	mem[12'h6CA] = 12'hF00;
	mem[12'h6CB] = 12'hF00;
	mem[12'h6CC] = 12'hF00;
	mem[12'h6CD] = 12'hF00;
	mem[12'h6CE] = 12'hF00;
	mem[12'h6CF] = 12'hF00;
	mem[12'h6D0] = 12'hF00;
	mem[12'h6D1] = 12'hF00;
	mem[12'h6D2] = 12'hF00;
	mem[12'h6D3] = 12'hF00;
	mem[12'h6D4] = 12'hFFF;
	mem[12'h6D5] = 12'hFFF;
	mem[12'h6D6] = 12'hFFF;
	mem[12'h6D7] = 12'hFFF;
	mem[12'h6D8] = 12'hFFF;
	mem[12'h6D9] = 12'hFFF;
	mem[12'h6DA] = 12'h01C;
	mem[12'h6DB] = 12'h00C;
	mem[12'h6DC] = 12'h00C;
	mem[12'h6DD] = 12'h00C;
	mem[12'h6DE] = 12'h00C;
	mem[12'h6DF] = 12'h01C;
	mem[12'h6E0] = 12'h01C;
	mem[12'h6E1] = 12'hE22;
	mem[12'h6E2] = 12'hF00;
	mem[12'h6E3] = 12'hF00;
	mem[12'h6E4] = 12'hF00;
	mem[12'h6E5] = 12'hF00;
	mem[12'h6E6] = 12'hF00;
	mem[12'h6E7] = 12'hF00;
	mem[12'h6E8] = 12'hF00;
	mem[12'h6E9] = 12'hFFF;
	mem[12'h6EA] = 12'hFFF;
	mem[12'h6EB] = 12'hFFF;
	mem[12'h6EC] = 12'hFFF;
	mem[12'h6ED] = 12'hFFF;
	mem[12'h6EE] = 12'h01C;
	mem[12'h6EF] = 12'h01C;
	mem[12'h6F0] = 12'h00C;
	mem[12'h6F1] = 12'h00C;
	mem[12'h6F2] = 12'h00C;
	mem[12'h6F3] = 12'h00C;
	mem[12'h6F4] = 12'h01C;
	mem[12'h6F5] = 12'hFFF;
	mem[12'h6F6] = 12'hF00;
	mem[12'h6F7] = 12'hF00;
	mem[12'h6F8] = 12'hE22;
	mem[12'h6F9] = 12'hFFF;
	mem[12'h6FA] = 12'hFFF;
	mem[12'h6FB] = 12'hFFF;
	mem[12'h6FC] = 12'hFFF;
	mem[12'h6FD] = 12'hFFF;
	mem[12'h6FE] = 12'hFFF;
	mem[12'h6FF] = 12'hFFF;
	mem[12'h700] = 12'hFFF;
	mem[12'h701] = 12'hFFF;
	mem[12'h702] = 12'hFFF;
	mem[12'h703] = 12'hFFF;
	mem[12'h704] = 12'hFFF;
	mem[12'h705] = 12'hFFF;
	mem[12'h706] = 12'hFFF;
	mem[12'h707] = 12'hE22;
	mem[12'h708] = 12'hF00;
	mem[12'h709] = 12'hF00;
	mem[12'h70A] = 12'hF00;
	mem[12'h70B] = 12'hF00;
	mem[12'h70C] = 12'hF00;
	mem[12'h70D] = 12'hF00;
	mem[12'h70E] = 12'hF00;
	mem[12'h70F] = 12'hF00;
	mem[12'h710] = 12'hF00;
	mem[12'h711] = 12'hF00;
	mem[12'h712] = 12'hF00;
	mem[12'h713] = 12'hF00;
	mem[12'h714] = 12'hFFF;
	mem[12'h715] = 12'hFFF;
	mem[12'h716] = 12'hFFF;
	mem[12'h717] = 12'hFFF;
	mem[12'h718] = 12'hFFF;
	mem[12'h719] = 12'hFFF;
	mem[12'h71A] = 12'h01C;
	mem[12'h71B] = 12'h01C;
	mem[12'h71C] = 12'h00C;
	mem[12'h71D] = 12'h00C;
	mem[12'h71E] = 12'h01C;
	mem[12'h71F] = 12'h01C;
	mem[12'h720] = 12'hFFF;
	mem[12'h721] = 12'hE22;
	mem[12'h722] = 12'hF00;
	mem[12'h723] = 12'hF00;
	mem[12'h724] = 12'hF00;
	mem[12'h725] = 12'hF00;
	mem[12'h726] = 12'hF00;
	mem[12'h727] = 12'hF00;
	mem[12'h728] = 12'hF00;
	mem[12'h729] = 12'hFFF;
	mem[12'h72A] = 12'hFFF;
	mem[12'h72B] = 12'hFFF;
	mem[12'h72C] = 12'hFFF;
	mem[12'h72D] = 12'hFFF;
	mem[12'h72E] = 12'hFFF;
	mem[12'h72F] = 12'h01C;
	mem[12'h730] = 12'h01C;
	mem[12'h731] = 12'h00C;
	mem[12'h732] = 12'h00C;
	mem[12'h733] = 12'h01C;
	mem[12'h734] = 12'h01C;
	mem[12'h735] = 12'hF00;
	mem[12'h736] = 12'hF00;
	mem[12'h737] = 12'hF00;
	mem[12'h738] = 12'hE22;
	mem[12'h739] = 12'hFFF;
	mem[12'h73A] = 12'hFFF;
	mem[12'h73B] = 12'hFFF;
	mem[12'h73C] = 12'hFFF;
	mem[12'h73D] = 12'hFFF;
	mem[12'h73E] = 12'hFFF;
	mem[12'h73F] = 12'hFFF;
	mem[12'h740] = 12'hFFF;
	mem[12'h741] = 12'hFFF;
	mem[12'h742] = 12'hFFF;
	mem[12'h743] = 12'hFFF;
	mem[12'h744] = 12'hFFF;
	mem[12'h745] = 12'hFFF;
	mem[12'h746] = 12'hFFF;
	mem[12'h747] = 12'hE22;
	mem[12'h748] = 12'hF00;
	mem[12'h749] = 12'hF00;
	mem[12'h74A] = 12'hF00;
	mem[12'h74B] = 12'hF00;
	mem[12'h74C] = 12'hF00;
	mem[12'h74D] = 12'hF00;
	mem[12'h74E] = 12'hF00;
	mem[12'h74F] = 12'hF00;
	mem[12'h750] = 12'hF00;
	mem[12'h751] = 12'hF00;
	mem[12'h752] = 12'hF00;
	mem[12'h753] = 12'hF00;
	mem[12'h754] = 12'hF00;
	mem[12'h755] = 12'hFFF;
	mem[12'h756] = 12'hFFF;
	mem[12'h757] = 12'hFFF;
	mem[12'h758] = 12'hFFF;
	mem[12'h759] = 12'hFFF;
	mem[12'h75A] = 12'hFFF;
	mem[12'h75B] = 12'h01C;
	mem[12'h75C] = 12'h01C;
	mem[12'h75D] = 12'h01C;
	mem[12'h75E] = 12'h01C;
	mem[12'h75F] = 12'hFFF;
	mem[12'h760] = 12'hF00;
	mem[12'h761] = 12'hF00;
	mem[12'h762] = 12'hF00;
	mem[12'h763] = 12'hF00;
	mem[12'h764] = 12'hF00;
	mem[12'h765] = 12'hF00;
	mem[12'h766] = 12'hF00;
	mem[12'h767] = 12'hF00;
	mem[12'h768] = 12'hE22;
	mem[12'h769] = 12'hFFF;
	mem[12'h76A] = 12'hFFF;
	mem[12'h76B] = 12'hFFF;
	mem[12'h76C] = 12'hFFF;
	mem[12'h76D] = 12'hFFF;
	mem[12'h76E] = 12'hFFF;
	mem[12'h76F] = 12'hFFF;
	mem[12'h770] = 12'h01C;
	mem[12'h771] = 12'h01C;
	mem[12'h772] = 12'h01C;
	mem[12'h773] = 12'h01C;
	mem[12'h774] = 12'hFFF;
	mem[12'h775] = 12'hE22;
	mem[12'h776] = 12'hF00;
	mem[12'h777] = 12'hF00;
	mem[12'h778] = 12'hE22;
	mem[12'h779] = 12'hFFF;
	mem[12'h77A] = 12'hFFF;
	mem[12'h77B] = 12'hFFF;
	mem[12'h77C] = 12'hFFF;
	mem[12'h77D] = 12'hFFF;
	mem[12'h77E] = 12'hFFF;
	mem[12'h77F] = 12'hFFF;
	mem[12'h780] = 12'hFFF;
	mem[12'h781] = 12'hFFF;
	mem[12'h782] = 12'hFFF;
	mem[12'h783] = 12'hFFF;
	mem[12'h784] = 12'hFFF;
	mem[12'h785] = 12'hFFF;
	mem[12'h786] = 12'hFFF;
	mem[12'h787] = 12'hE22;
	mem[12'h788] = 12'hF00;
	mem[12'h789] = 12'hF00;
	mem[12'h78A] = 12'hF00;
	mem[12'h78B] = 12'hF00;
	mem[12'h78C] = 12'hF00;
	mem[12'h78D] = 12'hF00;
	mem[12'h78E] = 12'hF00;
	mem[12'h78F] = 12'hF00;
	mem[12'h790] = 12'hF00;
	mem[12'h791] = 12'hF00;
	mem[12'h792] = 12'hF00;
	mem[12'h793] = 12'hF00;
	mem[12'h794] = 12'hF00;
	mem[12'h795] = 12'hFFF;
	mem[12'h796] = 12'hFFF;
	mem[12'h797] = 12'hFFF;
	mem[12'h798] = 12'hFFF;
	mem[12'h799] = 12'hFFF;
	mem[12'h79A] = 12'hFFF;
	mem[12'h79B] = 12'hFFF;
	mem[12'h79C] = 12'hFFF;
	mem[12'h79D] = 12'hFFF;
	mem[12'h79E] = 12'hFFF;
	mem[12'h79F] = 12'hFFF;
	mem[12'h7A0] = 12'hE22;
	mem[12'h7A1] = 12'hF00;
	mem[12'h7A2] = 12'hF00;
	mem[12'h7A3] = 12'hF00;
	mem[12'h7A4] = 12'hF00;
	mem[12'h7A5] = 12'hF00;
	mem[12'h7A6] = 12'hF00;
	mem[12'h7A7] = 12'hF00;
	mem[12'h7A8] = 12'hF00;
	mem[12'h7A9] = 12'hF00;
	mem[12'h7AA] = 12'hFFF;
	mem[12'h7AB] = 12'hFFF;
	mem[12'h7AC] = 12'hFFF;
	mem[12'h7AD] = 12'hFFF;
	mem[12'h7AE] = 12'hFFF;
	mem[12'h7AF] = 12'hFFF;
	mem[12'h7B0] = 12'hFFF;
	mem[12'h7B1] = 12'hFFF;
	mem[12'h7B2] = 12'hFFF;
	mem[12'h7B3] = 12'hFFF;
	mem[12'h7B4] = 12'hF00;
	mem[12'h7B5] = 12'hF00;
	mem[12'h7B6] = 12'hF00;
	mem[12'h7B7] = 12'hF00;
	mem[12'h7B8] = 12'hE22;
	mem[12'h7B9] = 12'hFFF;
	mem[12'h7BA] = 12'hFFF;
	mem[12'h7BB] = 12'hFFF;
	mem[12'h7BC] = 12'hFFF;
	mem[12'h7BD] = 12'hFFF;
	mem[12'h7BE] = 12'hFFF;
	mem[12'h7BF] = 12'hFFF;
	mem[12'h7C0] = 12'hFFF;
	mem[12'h7C1] = 12'hFFF;
	mem[12'h7C2] = 12'hFFF;
	mem[12'h7C3] = 12'hFFF;
	mem[12'h7C4] = 12'hFFF;
	mem[12'h7C5] = 12'hFFF;
	mem[12'h7C6] = 12'hFFF;
	mem[12'h7C7] = 12'hE22;
	mem[12'h7C8] = 12'hF00;
	mem[12'h7C9] = 12'hF00;
	mem[12'h7CA] = 12'hF00;
	mem[12'h7CB] = 12'hF00;
	mem[12'h7CC] = 12'hF00;
	mem[12'h7CD] = 12'hF00;
	mem[12'h7CE] = 12'hF00;
	mem[12'h7CF] = 12'hF00;
	mem[12'h7D0] = 12'hF00;
	mem[12'h7D1] = 12'hF00;
	mem[12'h7D2] = 12'hF00;
	mem[12'h7D3] = 12'hF00;
	mem[12'h7D4] = 12'hF00;
	mem[12'h7D5] = 12'hE22;
	mem[12'h7D6] = 12'hFFF;
	mem[12'h7D7] = 12'hFFF;
	mem[12'h7D8] = 12'hFFF;
	mem[12'h7D9] = 12'hFFF;
	mem[12'h7DA] = 12'hFFF;
	mem[12'h7DB] = 12'hFFF;
	mem[12'h7DC] = 12'hFFF;
	mem[12'h7DD] = 12'hFFF;
	mem[12'h7DE] = 12'hFFF;
	mem[12'h7DF] = 12'hE22;
	mem[12'h7E0] = 12'hF00;
	mem[12'h7E1] = 12'hF00;
	mem[12'h7E2] = 12'hF00;
	mem[12'h7E3] = 12'hF00;
	mem[12'h7E4] = 12'hF00;
	mem[12'h7E5] = 12'hF00;
	mem[12'h7E6] = 12'hF00;
	mem[12'h7E7] = 12'hF00;
	mem[12'h7E8] = 12'hF00;
	mem[12'h7E9] = 12'hF00;
	mem[12'h7EA] = 12'hF00;
	mem[12'h7EB] = 12'hFFF;
	mem[12'h7EC] = 12'hFFF;
	mem[12'h7ED] = 12'hFFF;
	mem[12'h7EE] = 12'hFFF;
	mem[12'h7EF] = 12'hFFF;
	mem[12'h7F0] = 12'hFFF;
	mem[12'h7F1] = 12'hFFF;
	mem[12'h7F2] = 12'hFFF;
	mem[12'h7F3] = 12'hFFF;
	mem[12'h7F4] = 12'hF00;
	mem[12'h7F5] = 12'hF00;
	mem[12'h7F6] = 12'hF00;
	mem[12'h7F7] = 12'hF00;
	mem[12'h7F8] = 12'hE22;
	mem[12'h7F9] = 12'hFFF;
	mem[12'h7FA] = 12'hFFF;
	mem[12'h7FB] = 12'hFFF;
	mem[12'h7FC] = 12'hFFF;
	mem[12'h7FD] = 12'hFFF;
	mem[12'h7FE] = 12'hFFF;
	mem[12'h7FF] = 12'hFFF;
	mem[12'h800] = 12'hFFF;
	mem[12'h801] = 12'hFFF;
	mem[12'h802] = 12'hFFF;
	mem[12'h803] = 12'hFFF;
	mem[12'h804] = 12'hFFF;
	mem[12'h805] = 12'hFFF;
	mem[12'h806] = 12'hFFF;
	mem[12'h807] = 12'hE22;
	mem[12'h808] = 12'hF00;
	mem[12'h809] = 12'hF00;
	mem[12'h80A] = 12'hF00;
	mem[12'h80B] = 12'hF00;
	mem[12'h80C] = 12'hF00;
	mem[12'h80D] = 12'hF00;
	mem[12'h80E] = 12'hF00;
	mem[12'h80F] = 12'hF00;
	mem[12'h810] = 12'hF00;
	mem[12'h811] = 12'hF00;
	mem[12'h812] = 12'hF00;
	mem[12'h813] = 12'hF00;
	mem[12'h814] = 12'hF00;
	mem[12'h815] = 12'hF00;
	mem[12'h816] = 12'hE22;
	mem[12'h817] = 12'hF00;
	mem[12'h818] = 12'hFFF;
	mem[12'h819] = 12'hFFF;
	mem[12'h81A] = 12'hFFF;
	mem[12'h81B] = 12'hFFF;
	mem[12'h81C] = 12'hFFF;
	mem[12'h81D] = 12'hFFF;
	mem[12'h81E] = 12'hE22;
	mem[12'h81F] = 12'hF00;
	mem[12'h820] = 12'hF00;
	mem[12'h821] = 12'hF00;
	mem[12'h822] = 12'hF00;
	mem[12'h823] = 12'hF00;
	mem[12'h824] = 12'hF00;
	mem[12'h825] = 12'hF00;
	mem[12'h826] = 12'hF00;
	mem[12'h827] = 12'hF00;
	mem[12'h828] = 12'hF00;
	mem[12'h829] = 12'hF00;
	mem[12'h82A] = 12'hF00;
	mem[12'h82B] = 12'hF00;
	mem[12'h82C] = 12'hFFF;
	mem[12'h82D] = 12'hFFF;
	mem[12'h82E] = 12'hFFF;
	mem[12'h82F] = 12'hFFF;
	mem[12'h830] = 12'hFFF;
	mem[12'h831] = 12'hFFF;
	mem[12'h832] = 12'hF00;
	mem[12'h833] = 12'hF00;
	mem[12'h834] = 12'hF00;
	mem[12'h835] = 12'hF00;
	mem[12'h836] = 12'hF00;
	mem[12'h837] = 12'hF00;
	mem[12'h838] = 12'hE22;
	mem[12'h839] = 12'hFFF;
	mem[12'h83A] = 12'hFFF;
	mem[12'h83B] = 12'hFFF;
	mem[12'h83C] = 12'hFFF;
	mem[12'h83D] = 12'hFFF;
	mem[12'h83E] = 12'hFFF;
	mem[12'h83F] = 12'hFFF;
	mem[12'h840] = 12'hFFF;
	mem[12'h841] = 12'hFFF;
	mem[12'h842] = 12'hFFF;
	mem[12'h843] = 12'hFFF;
	mem[12'h844] = 12'hFFF;
	mem[12'h845] = 12'hFFF;
	mem[12'h846] = 12'hFFF;
	mem[12'h847] = 12'hE22;
	mem[12'h848] = 12'hF00;
	mem[12'h849] = 12'hF00;
	mem[12'h84A] = 12'hF00;
	mem[12'h84B] = 12'hF00;
	mem[12'h84C] = 12'hF00;
	mem[12'h84D] = 12'hF00;
	mem[12'h84E] = 12'hF00;
	mem[12'h84F] = 12'hF00;
	mem[12'h850] = 12'hF00;
	mem[12'h851] = 12'hF00;
	mem[12'h852] = 12'hF00;
	mem[12'h853] = 12'hF00;
	mem[12'h854] = 12'hF00;
	mem[12'h855] = 12'hF00;
	mem[12'h856] = 12'hF00;
	mem[12'h857] = 12'hF00;
	mem[12'h858] = 12'hE22;
	mem[12'h859] = 12'hE22;
	mem[12'h85A] = 12'hF00;
	mem[12'h85B] = 12'hF00;
	mem[12'h85C] = 12'hE22;
	mem[12'h85D] = 12'hF00;
	mem[12'h85E] = 12'hF00;
	mem[12'h85F] = 12'hF00;
	mem[12'h860] = 12'hF00;
	mem[12'h861] = 12'hF00;
	mem[12'h862] = 12'hF00;
	mem[12'h863] = 12'hF00;
	mem[12'h864] = 12'hF00;
	mem[12'h865] = 12'hF00;
	mem[12'h866] = 12'hF00;
	mem[12'h867] = 12'hF00;
	mem[12'h868] = 12'hF00;
	mem[12'h869] = 12'hF00;
	mem[12'h86A] = 12'hF00;
	mem[12'h86B] = 12'hF00;
	mem[12'h86C] = 12'hF00;
	mem[12'h86D] = 12'hE22;
	mem[12'h86E] = 12'hF00;
	mem[12'h86F] = 12'hF00;
	mem[12'h870] = 12'hE22;
	mem[12'h871] = 12'hE22;
	mem[12'h872] = 12'hF00;
	mem[12'h873] = 12'hF00;
	mem[12'h874] = 12'hF00;
	mem[12'h875] = 12'hF00;
	mem[12'h876] = 12'hF00;
	mem[12'h877] = 12'hF00;
	mem[12'h878] = 12'hE22;
	mem[12'h879] = 12'hFFF;
	mem[12'h87A] = 12'hFFF;
	mem[12'h87B] = 12'hFFF;
	mem[12'h87C] = 12'hFFF;
	mem[12'h87D] = 12'hFFF;
	mem[12'h87E] = 12'hFFF;
	mem[12'h87F] = 12'hFFF;
	mem[12'h880] = 12'hFFF;
	mem[12'h881] = 12'hFFF;
	mem[12'h882] = 12'hFFF;
	mem[12'h883] = 12'hFFF;
	mem[12'h884] = 12'hFFF;
	mem[12'h885] = 12'hFFF;
	mem[12'h886] = 12'hFFF;
	mem[12'h887] = 12'hE22;
	mem[12'h888] = 12'hF00;
	mem[12'h889] = 12'hF00;
	mem[12'h88A] = 12'hF00;
	mem[12'h88B] = 12'hF00;
	mem[12'h88C] = 12'hF00;
	mem[12'h88D] = 12'hF00;
	mem[12'h88E] = 12'hF00;
	mem[12'h88F] = 12'hF00;
	mem[12'h890] = 12'hF00;
	mem[12'h891] = 12'hF00;
	mem[12'h892] = 12'hF00;
	mem[12'h893] = 12'hF00;
	mem[12'h894] = 12'hF00;
	mem[12'h895] = 12'hF00;
	mem[12'h896] = 12'hF00;
	mem[12'h897] = 12'hF00;
	mem[12'h898] = 12'hF00;
	mem[12'h899] = 12'hF00;
	mem[12'h89A] = 12'hF00;
	mem[12'h89B] = 12'hF00;
	mem[12'h89C] = 12'hF00;
	mem[12'h89D] = 12'hF00;
	mem[12'h89E] = 12'hF00;
	mem[12'h89F] = 12'hF00;
	mem[12'h8A0] = 12'hF00;
	mem[12'h8A1] = 12'hF00;
	mem[12'h8A2] = 12'hF00;
	mem[12'h8A3] = 12'hF00;
	mem[12'h8A4] = 12'hF00;
	mem[12'h8A5] = 12'hF00;
	mem[12'h8A6] = 12'hF00;
	mem[12'h8A7] = 12'hF00;
	mem[12'h8A8] = 12'hF00;
	mem[12'h8A9] = 12'hF00;
	mem[12'h8AA] = 12'hF00;
	mem[12'h8AB] = 12'hF00;
	mem[12'h8AC] = 12'hF00;
	mem[12'h8AD] = 12'hF00;
	mem[12'h8AE] = 12'hF00;
	mem[12'h8AF] = 12'hF00;
	mem[12'h8B0] = 12'hF00;
	mem[12'h8B1] = 12'hF00;
	mem[12'h8B2] = 12'hF00;
	mem[12'h8B3] = 12'hF00;
	mem[12'h8B4] = 12'hF00;
	mem[12'h8B5] = 12'hF00;
	mem[12'h8B6] = 12'hF00;
	mem[12'h8B7] = 12'hF00;
	mem[12'h8B8] = 12'hE22;
	mem[12'h8B9] = 12'hFFF;
	mem[12'h8BA] = 12'hFFF;
	mem[12'h8BB] = 12'hFFF;
	mem[12'h8BC] = 12'hFFF;
	mem[12'h8BD] = 12'hFFF;
	mem[12'h8BE] = 12'hFFF;
	mem[12'h8BF] = 12'hFFF;
	mem[12'h8C0] = 12'hFFF;
	mem[12'h8C1] = 12'hFFF;
	mem[12'h8C2] = 12'hFFF;
	mem[12'h8C3] = 12'hFFF;
	mem[12'h8C4] = 12'hFFF;
	mem[12'h8C5] = 12'hFFF;
	mem[12'h8C6] = 12'hFFF;
	mem[12'h8C7] = 12'hE22;
	mem[12'h8C8] = 12'hF00;
	mem[12'h8C9] = 12'hF00;
	mem[12'h8CA] = 12'hF00;
	mem[12'h8CB] = 12'hF00;
	mem[12'h8CC] = 12'hF00;
	mem[12'h8CD] = 12'hF00;
	mem[12'h8CE] = 12'hF00;
	mem[12'h8CF] = 12'hF00;
	mem[12'h8D0] = 12'hF00;
	mem[12'h8D1] = 12'hF00;
	mem[12'h8D2] = 12'hF00;
	mem[12'h8D3] = 12'hF00;
	mem[12'h8D4] = 12'hF00;
	mem[12'h8D5] = 12'hF00;
	mem[12'h8D6] = 12'hF00;
	mem[12'h8D7] = 12'hF00;
	mem[12'h8D8] = 12'hF00;
	mem[12'h8D9] = 12'hF00;
	mem[12'h8DA] = 12'hF00;
	mem[12'h8DB] = 12'hF00;
	mem[12'h8DC] = 12'hF00;
	mem[12'h8DD] = 12'hF00;
	mem[12'h8DE] = 12'hF00;
	mem[12'h8DF] = 12'hF00;
	mem[12'h8E0] = 12'hF00;
	mem[12'h8E1] = 12'hF00;
	mem[12'h8E2] = 12'hF00;
	mem[12'h8E3] = 12'hF00;
	mem[12'h8E4] = 12'hF00;
	mem[12'h8E5] = 12'hF00;
	mem[12'h8E6] = 12'hF00;
	mem[12'h8E7] = 12'hF00;
	mem[12'h8E8] = 12'hF00;
	mem[12'h8E9] = 12'hF00;
	mem[12'h8EA] = 12'hF00;
	mem[12'h8EB] = 12'hF00;
	mem[12'h8EC] = 12'hF00;
	mem[12'h8ED] = 12'hF00;
	mem[12'h8EE] = 12'hF00;
	mem[12'h8EF] = 12'hF00;
	mem[12'h8F0] = 12'hF00;
	mem[12'h8F1] = 12'hF00;
	mem[12'h8F2] = 12'hF00;
	mem[12'h8F3] = 12'hF00;
	mem[12'h8F4] = 12'hF00;
	mem[12'h8F5] = 12'hF00;
	mem[12'h8F6] = 12'hF00;
	mem[12'h8F7] = 12'hF00;
	mem[12'h8F8] = 12'hE22;
	mem[12'h8F9] = 12'hFFF;
	mem[12'h8FA] = 12'hFFF;
	mem[12'h8FB] = 12'hFFF;
	mem[12'h8FC] = 12'hFFF;
	mem[12'h8FD] = 12'hFFF;
	mem[12'h8FE] = 12'hFFF;
	mem[12'h8FF] = 12'hFFF;
	mem[12'h900] = 12'hFFF;
	mem[12'h901] = 12'hFFF;
	mem[12'h902] = 12'hFFF;
	mem[12'h903] = 12'hFFF;
	mem[12'h904] = 12'hFFF;
	mem[12'h905] = 12'hFFF;
	mem[12'h906] = 12'hFFF;
	mem[12'h907] = 12'hE22;
	mem[12'h908] = 12'hF00;
	mem[12'h909] = 12'hF00;
	mem[12'h90A] = 12'hF00;
	mem[12'h90B] = 12'hF00;
	mem[12'h90C] = 12'hF00;
	mem[12'h90D] = 12'hF00;
	mem[12'h90E] = 12'hF00;
	mem[12'h90F] = 12'hF00;
	mem[12'h910] = 12'hF00;
	mem[12'h911] = 12'hF00;
	mem[12'h912] = 12'hF00;
	mem[12'h913] = 12'hF00;
	mem[12'h914] = 12'hF00;
	mem[12'h915] = 12'hF00;
	mem[12'h916] = 12'hF00;
	mem[12'h917] = 12'hF00;
	mem[12'h918] = 12'hF00;
	mem[12'h919] = 12'hF00;
	mem[12'h91A] = 12'hF00;
	mem[12'h91B] = 12'hF00;
	mem[12'h91C] = 12'hF00;
	mem[12'h91D] = 12'hF00;
	mem[12'h91E] = 12'hF00;
	mem[12'h91F] = 12'hF00;
	mem[12'h920] = 12'hF00;
	mem[12'h921] = 12'hF00;
	mem[12'h922] = 12'hF00;
	mem[12'h923] = 12'hF00;
	mem[12'h924] = 12'hF00;
	mem[12'h925] = 12'hF00;
	mem[12'h926] = 12'hF00;
	mem[12'h927] = 12'hF00;
	mem[12'h928] = 12'hF00;
	mem[12'h929] = 12'hF00;
	mem[12'h92A] = 12'hF00;
	mem[12'h92B] = 12'hF00;
	mem[12'h92C] = 12'hF00;
	mem[12'h92D] = 12'hF00;
	mem[12'h92E] = 12'hF00;
	mem[12'h92F] = 12'hF00;
	mem[12'h930] = 12'hF00;
	mem[12'h931] = 12'hF00;
	mem[12'h932] = 12'hF00;
	mem[12'h933] = 12'hF00;
	mem[12'h934] = 12'hF00;
	mem[12'h935] = 12'hF00;
	mem[12'h936] = 12'hF00;
	mem[12'h937] = 12'hF00;
	mem[12'h938] = 12'hE22;
	mem[12'h939] = 12'hFFF;
	mem[12'h93A] = 12'hFFF;
	mem[12'h93B] = 12'hFFF;
	mem[12'h93C] = 12'hFFF;
	mem[12'h93D] = 12'hFFF;
	mem[12'h93E] = 12'hFFF;
	mem[12'h93F] = 12'hFFF;
	mem[12'h940] = 12'hFFF;
	mem[12'h941] = 12'hFFF;
	mem[12'h942] = 12'hFFF;
	mem[12'h943] = 12'hFFF;
	mem[12'h944] = 12'hFFF;
	mem[12'h945] = 12'hFFF;
	mem[12'h946] = 12'hFFF;
	mem[12'h947] = 12'hE22;
	mem[12'h948] = 12'hF00;
	mem[12'h949] = 12'hF00;
	mem[12'h94A] = 12'hF00;
	mem[12'h94B] = 12'hF00;
	mem[12'h94C] = 12'hF00;
	mem[12'h94D] = 12'hF00;
	mem[12'h94E] = 12'hF00;
	mem[12'h94F] = 12'hF00;
	mem[12'h950] = 12'hF00;
	mem[12'h951] = 12'hF00;
	mem[12'h952] = 12'hF00;
	mem[12'h953] = 12'hF00;
	mem[12'h954] = 12'hF00;
	mem[12'h955] = 12'hF00;
	mem[12'h956] = 12'hF00;
	mem[12'h957] = 12'hF00;
	mem[12'h958] = 12'hF00;
	mem[12'h959] = 12'hF00;
	mem[12'h95A] = 12'hF00;
	mem[12'h95B] = 12'hF00;
	mem[12'h95C] = 12'hF00;
	mem[12'h95D] = 12'hF00;
	mem[12'h95E] = 12'hF00;
	mem[12'h95F] = 12'hF00;
	mem[12'h960] = 12'hF00;
	mem[12'h961] = 12'hF00;
	mem[12'h962] = 12'hF00;
	mem[12'h963] = 12'hF00;
	mem[12'h964] = 12'hF00;
	mem[12'h965] = 12'hF00;
	mem[12'h966] = 12'hF00;
	mem[12'h967] = 12'hF00;
	mem[12'h968] = 12'hF00;
	mem[12'h969] = 12'hF00;
	mem[12'h96A] = 12'hF00;
	mem[12'h96B] = 12'hF00;
	mem[12'h96C] = 12'hF00;
	mem[12'h96D] = 12'hF00;
	mem[12'h96E] = 12'hF00;
	mem[12'h96F] = 12'hF00;
	mem[12'h970] = 12'hF00;
	mem[12'h971] = 12'hF00;
	mem[12'h972] = 12'hF00;
	mem[12'h973] = 12'hF00;
	mem[12'h974] = 12'hF00;
	mem[12'h975] = 12'hF00;
	mem[12'h976] = 12'hF00;
	mem[12'h977] = 12'hF00;
	mem[12'h978] = 12'hE22;
	mem[12'h979] = 12'hFFF;
	mem[12'h97A] = 12'hFFF;
	mem[12'h97B] = 12'hFFF;
	mem[12'h97C] = 12'hFFF;
	mem[12'h97D] = 12'hFFF;
	mem[12'h97E] = 12'hFFF;
	mem[12'h97F] = 12'hFFF;
	mem[12'h980] = 12'hFFF;
	mem[12'h981] = 12'hFFF;
	mem[12'h982] = 12'hFFF;
	mem[12'h983] = 12'hFFF;
	mem[12'h984] = 12'hFFF;
	mem[12'h985] = 12'hFFF;
	mem[12'h986] = 12'hFFF;
	mem[12'h987] = 12'hE22;
	mem[12'h988] = 12'hF00;
	mem[12'h989] = 12'hF00;
	mem[12'h98A] = 12'hF00;
	mem[12'h98B] = 12'hF00;
	mem[12'h98C] = 12'hF00;
	mem[12'h98D] = 12'hF00;
	mem[12'h98E] = 12'hF00;
	mem[12'h98F] = 12'hF00;
	mem[12'h990] = 12'hF00;
	mem[12'h991] = 12'hF00;
	mem[12'h992] = 12'hF00;
	mem[12'h993] = 12'hF00;
	mem[12'h994] = 12'hF00;
	mem[12'h995] = 12'hF00;
	mem[12'h996] = 12'hF00;
	mem[12'h997] = 12'hF00;
	mem[12'h998] = 12'hF00;
	mem[12'h999] = 12'hF00;
	mem[12'h99A] = 12'hF00;
	mem[12'h99B] = 12'hF00;
	mem[12'h99C] = 12'hF00;
	mem[12'h99D] = 12'hF00;
	mem[12'h99E] = 12'hF00;
	mem[12'h99F] = 12'hF00;
	mem[12'h9A0] = 12'hF00;
	mem[12'h9A1] = 12'hF00;
	mem[12'h9A2] = 12'hF00;
	mem[12'h9A3] = 12'hF00;
	mem[12'h9A4] = 12'hF00;
	mem[12'h9A5] = 12'hF00;
	mem[12'h9A6] = 12'hF00;
	mem[12'h9A7] = 12'hF00;
	mem[12'h9A8] = 12'hF00;
	mem[12'h9A9] = 12'hF00;
	mem[12'h9AA] = 12'hF00;
	mem[12'h9AB] = 12'hF00;
	mem[12'h9AC] = 12'hF00;
	mem[12'h9AD] = 12'hF00;
	mem[12'h9AE] = 12'hF00;
	mem[12'h9AF] = 12'hF00;
	mem[12'h9B0] = 12'hF00;
	mem[12'h9B1] = 12'hF00;
	mem[12'h9B2] = 12'hF00;
	mem[12'h9B3] = 12'hF00;
	mem[12'h9B4] = 12'hF00;
	mem[12'h9B5] = 12'hF00;
	mem[12'h9B6] = 12'hF00;
	mem[12'h9B7] = 12'hF00;
	mem[12'h9B8] = 12'hE22;
	mem[12'h9B9] = 12'hFFF;
	mem[12'h9BA] = 12'hFFF;
	mem[12'h9BB] = 12'hFFF;
	mem[12'h9BC] = 12'hFFF;
	mem[12'h9BD] = 12'hFFF;
	mem[12'h9BE] = 12'hFFF;
	mem[12'h9BF] = 12'hFFF;
	mem[12'h9C0] = 12'hFFF;
	mem[12'h9C1] = 12'hFFF;
	mem[12'h9C2] = 12'hFFF;
	mem[12'h9C3] = 12'hFFF;
	mem[12'h9C4] = 12'hFFF;
	mem[12'h9C5] = 12'hFFF;
	mem[12'h9C6] = 12'hFFF;
	mem[12'h9C7] = 12'hE22;
	mem[12'h9C8] = 12'hF00;
	mem[12'h9C9] = 12'hF00;
	mem[12'h9CA] = 12'hF00;
	mem[12'h9CB] = 12'hF00;
	mem[12'h9CC] = 12'hF00;
	mem[12'h9CD] = 12'hF00;
	mem[12'h9CE] = 12'hF00;
	mem[12'h9CF] = 12'hF00;
	mem[12'h9D0] = 12'hF00;
	mem[12'h9D1] = 12'hF00;
	mem[12'h9D2] = 12'hF00;
	mem[12'h9D3] = 12'hF00;
	mem[12'h9D4] = 12'hF00;
	mem[12'h9D5] = 12'hF00;
	mem[12'h9D6] = 12'hF00;
	mem[12'h9D7] = 12'hF00;
	mem[12'h9D8] = 12'hF00;
	mem[12'h9D9] = 12'hF00;
	mem[12'h9DA] = 12'hF00;
	mem[12'h9DB] = 12'hF00;
	mem[12'h9DC] = 12'hF00;
	mem[12'h9DD] = 12'hF00;
	mem[12'h9DE] = 12'hF00;
	mem[12'h9DF] = 12'hF00;
	mem[12'h9E0] = 12'hF00;
	mem[12'h9E1] = 12'hF00;
	mem[12'h9E2] = 12'hF00;
	mem[12'h9E3] = 12'hF00;
	mem[12'h9E4] = 12'hF00;
	mem[12'h9E5] = 12'hF00;
	mem[12'h9E6] = 12'hF00;
	mem[12'h9E7] = 12'hF00;
	mem[12'h9E8] = 12'hF00;
	mem[12'h9E9] = 12'hF00;
	mem[12'h9EA] = 12'hF00;
	mem[12'h9EB] = 12'hF00;
	mem[12'h9EC] = 12'hF00;
	mem[12'h9ED] = 12'hF00;
	mem[12'h9EE] = 12'hF00;
	mem[12'h9EF] = 12'hF00;
	mem[12'h9F0] = 12'hF00;
	mem[12'h9F1] = 12'hF00;
	mem[12'h9F2] = 12'hF00;
	mem[12'h9F3] = 12'hF00;
	mem[12'h9F4] = 12'hF00;
	mem[12'h9F5] = 12'hF00;
	mem[12'h9F6] = 12'hF00;
	mem[12'h9F7] = 12'hF00;
	mem[12'h9F8] = 12'hE22;
	mem[12'h9F9] = 12'hFFF;
	mem[12'h9FA] = 12'hFFF;
	mem[12'h9FB] = 12'hFFF;
	mem[12'h9FC] = 12'hFFF;
	mem[12'h9FD] = 12'hFFF;
	mem[12'h9FE] = 12'hFFF;
	mem[12'h9FF] = 12'hFFF;
	mem[12'hA00] = 12'hFFF;
	mem[12'hA01] = 12'hFFF;
	mem[12'hA02] = 12'hFFF;
	mem[12'hA03] = 12'hFFF;
	mem[12'hA04] = 12'hFFF;
	mem[12'hA05] = 12'hFFF;
	mem[12'hA06] = 12'hFFF;
	mem[12'hA07] = 12'hE22;
	mem[12'hA08] = 12'hF00;
	mem[12'hA09] = 12'hF00;
	mem[12'hA0A] = 12'hF00;
	mem[12'hA0B] = 12'hF00;
	mem[12'hA0C] = 12'hF00;
	mem[12'hA0D] = 12'hF00;
	mem[12'hA0E] = 12'hF00;
	mem[12'hA0F] = 12'hF00;
	mem[12'hA10] = 12'hF00;
	mem[12'hA11] = 12'hF00;
	mem[12'hA12] = 12'hF00;
	mem[12'hA13] = 12'hF00;
	mem[12'hA14] = 12'hF00;
	mem[12'hA15] = 12'hF00;
	mem[12'hA16] = 12'hF00;
	mem[12'hA17] = 12'hF00;
	mem[12'hA18] = 12'hF00;
	mem[12'hA19] = 12'hF00;
	mem[12'hA1A] = 12'hF00;
	mem[12'hA1B] = 12'hF00;
	mem[12'hA1C] = 12'hF00;
	mem[12'hA1D] = 12'hF00;
	mem[12'hA1E] = 12'hF00;
	mem[12'hA1F] = 12'hF00;
	mem[12'hA20] = 12'hF00;
	mem[12'hA21] = 12'hF00;
	mem[12'hA22] = 12'hF00;
	mem[12'hA23] = 12'hF00;
	mem[12'hA24] = 12'hF00;
	mem[12'hA25] = 12'hF00;
	mem[12'hA26] = 12'hF00;
	mem[12'hA27] = 12'hF00;
	mem[12'hA28] = 12'hF00;
	mem[12'hA29] = 12'hF00;
	mem[12'hA2A] = 12'hF00;
	mem[12'hA2B] = 12'hF00;
	mem[12'hA2C] = 12'hF00;
	mem[12'hA2D] = 12'hF00;
	mem[12'hA2E] = 12'hF00;
	mem[12'hA2F] = 12'hF00;
	mem[12'hA30] = 12'hF00;
	mem[12'hA31] = 12'hF00;
	mem[12'hA32] = 12'hF00;
	mem[12'hA33] = 12'hF00;
	mem[12'hA34] = 12'hF00;
	mem[12'hA35] = 12'hF00;
	mem[12'hA36] = 12'hF00;
	mem[12'hA37] = 12'hF00;
	mem[12'hA38] = 12'hE22;
	mem[12'hA39] = 12'hFFF;
	mem[12'hA3A] = 12'hFFF;
	mem[12'hA3B] = 12'hFFF;
	mem[12'hA3C] = 12'hFFF;
	mem[12'hA3D] = 12'hFFF;
	mem[12'hA3E] = 12'hFFF;
	mem[12'hA3F] = 12'hFFF;
	mem[12'hA40] = 12'hFFF;
	mem[12'hA41] = 12'hFFF;
	mem[12'hA42] = 12'hFFF;
	mem[12'hA43] = 12'hFFF;
	mem[12'hA44] = 12'hFFF;
	mem[12'hA45] = 12'hFFF;
	mem[12'hA46] = 12'hFFF;
	mem[12'hA47] = 12'hE22;
	mem[12'hA48] = 12'hF00;
	mem[12'hA49] = 12'hF00;
	mem[12'hA4A] = 12'hF00;
	mem[12'hA4B] = 12'hF00;
	mem[12'hA4C] = 12'hF00;
	mem[12'hA4D] = 12'hF00;
	mem[12'hA4E] = 12'hF00;
	mem[12'hA4F] = 12'hF00;
	mem[12'hA50] = 12'hF00;
	mem[12'hA51] = 12'hF00;
	mem[12'hA52] = 12'hF00;
	mem[12'hA53] = 12'hF00;
	mem[12'hA54] = 12'hF00;
	mem[12'hA55] = 12'hF00;
	mem[12'hA56] = 12'hF00;
	mem[12'hA57] = 12'hF00;
	mem[12'hA58] = 12'hF00;
	mem[12'hA59] = 12'hF00;
	mem[12'hA5A] = 12'hF00;
	mem[12'hA5B] = 12'hF00;
	mem[12'hA5C] = 12'hF00;
	mem[12'hA5D] = 12'hF00;
	mem[12'hA5E] = 12'hF00;
	mem[12'hA5F] = 12'hF00;
	mem[12'hA60] = 12'hF00;
	mem[12'hA61] = 12'hF00;
	mem[12'hA62] = 12'hF00;
	mem[12'hA63] = 12'hF00;
	mem[12'hA64] = 12'hF00;
	mem[12'hA65] = 12'hF00;
	mem[12'hA66] = 12'hF00;
	mem[12'hA67] = 12'hF00;
	mem[12'hA68] = 12'hF00;
	mem[12'hA69] = 12'hF00;
	mem[12'hA6A] = 12'hF00;
	mem[12'hA6B] = 12'hF00;
	mem[12'hA6C] = 12'hF00;
	mem[12'hA6D] = 12'hF00;
	mem[12'hA6E] = 12'hF00;
	mem[12'hA6F] = 12'hF00;
	mem[12'hA70] = 12'hF00;
	mem[12'hA71] = 12'hF00;
	mem[12'hA72] = 12'hF00;
	mem[12'hA73] = 12'hF00;
	mem[12'hA74] = 12'hF00;
	mem[12'hA75] = 12'hF00;
	mem[12'hA76] = 12'hF00;
	mem[12'hA77] = 12'hF00;
	mem[12'hA78] = 12'hE22;
	mem[12'hA79] = 12'hFFF;
	mem[12'hA7A] = 12'hFFF;
	mem[12'hA7B] = 12'hFFF;
	mem[12'hA7C] = 12'hFFF;
	mem[12'hA7D] = 12'hFFF;
	mem[12'hA7E] = 12'hFFF;
	mem[12'hA7F] = 12'hFFF;
	mem[12'hA80] = 12'hFFF;
	mem[12'hA81] = 12'hFFF;
	mem[12'hA82] = 12'hFFF;
	mem[12'hA83] = 12'hFFF;
	mem[12'hA84] = 12'hFFF;
	mem[12'hA85] = 12'hFFF;
	mem[12'hA86] = 12'hFFF;
	mem[12'hA87] = 12'hE22;
	mem[12'hA88] = 12'hF00;
	mem[12'hA89] = 12'hF00;
	mem[12'hA8A] = 12'hF00;
	mem[12'hA8B] = 12'hF00;
	mem[12'hA8C] = 12'hF00;
	mem[12'hA8D] = 12'hF00;
	mem[12'hA8E] = 12'hF00;
	mem[12'hA8F] = 12'hF00;
	mem[12'hA90] = 12'hF00;
	mem[12'hA91] = 12'hF00;
	mem[12'hA92] = 12'hF00;
	mem[12'hA93] = 12'hF00;
	mem[12'hA94] = 12'hF00;
	mem[12'hA95] = 12'hF00;
	mem[12'hA96] = 12'hF00;
	mem[12'hA97] = 12'hF00;
	mem[12'hA98] = 12'hF00;
	mem[12'hA99] = 12'hF00;
	mem[12'hA9A] = 12'hF00;
	mem[12'hA9B] = 12'hF00;
	mem[12'hA9C] = 12'hF00;
	mem[12'hA9D] = 12'hF00;
	mem[12'hA9E] = 12'hF00;
	mem[12'hA9F] = 12'hF00;
	mem[12'hAA0] = 12'hF00;
	mem[12'hAA1] = 12'hF00;
	mem[12'hAA2] = 12'hF00;
	mem[12'hAA3] = 12'hF00;
	mem[12'hAA4] = 12'hF00;
	mem[12'hAA5] = 12'hF00;
	mem[12'hAA6] = 12'hF00;
	mem[12'hAA7] = 12'hF00;
	mem[12'hAA8] = 12'hF00;
	mem[12'hAA9] = 12'hF00;
	mem[12'hAAA] = 12'hF00;
	mem[12'hAAB] = 12'hF00;
	mem[12'hAAC] = 12'hF00;
	mem[12'hAAD] = 12'hF00;
	mem[12'hAAE] = 12'hF00;
	mem[12'hAAF] = 12'hF00;
	mem[12'hAB0] = 12'hF00;
	mem[12'hAB1] = 12'hF00;
	mem[12'hAB2] = 12'hF00;
	mem[12'hAB3] = 12'hF00;
	mem[12'hAB4] = 12'hF00;
	mem[12'hAB5] = 12'hF00;
	mem[12'hAB6] = 12'hF00;
	mem[12'hAB7] = 12'hF00;
	mem[12'hAB8] = 12'hE22;
	mem[12'hAB9] = 12'hFFF;
	mem[12'hABA] = 12'hFFF;
	mem[12'hABB] = 12'hFFF;
	mem[12'hABC] = 12'hFFF;
	mem[12'hABD] = 12'hFFF;
	mem[12'hABE] = 12'hFFF;
	mem[12'hABF] = 12'hFFF;
	mem[12'hAC0] = 12'hFFF;
	mem[12'hAC1] = 12'hFFF;
	mem[12'hAC2] = 12'hFFF;
	mem[12'hAC3] = 12'hFFF;
	mem[12'hAC4] = 12'hFFF;
	mem[12'hAC5] = 12'hFFF;
	mem[12'hAC6] = 12'hFFF;
	mem[12'hAC7] = 12'hE22;
	mem[12'hAC8] = 12'hF00;
	mem[12'hAC9] = 12'hF00;
	mem[12'hACA] = 12'hF00;
	mem[12'hACB] = 12'hF00;
	mem[12'hACC] = 12'hF00;
	mem[12'hACD] = 12'hF00;
	mem[12'hACE] = 12'hF00;
	mem[12'hACF] = 12'hF00;
	mem[12'hAD0] = 12'hF00;
	mem[12'hAD1] = 12'hF00;
	mem[12'hAD2] = 12'hF00;
	mem[12'hAD3] = 12'hF00;
	mem[12'hAD4] = 12'hF00;
	mem[12'hAD5] = 12'hF00;
	mem[12'hAD6] = 12'hF00;
	mem[12'hAD7] = 12'hF00;
	mem[12'hAD8] = 12'hF00;
	mem[12'hAD9] = 12'hF00;
	mem[12'hADA] = 12'hF00;
	mem[12'hADB] = 12'hF00;
	mem[12'hADC] = 12'hF00;
	mem[12'hADD] = 12'hF00;
	mem[12'hADE] = 12'hF00;
	mem[12'hADF] = 12'hF00;
	mem[12'hAE0] = 12'hF00;
	mem[12'hAE1] = 12'hF00;
	mem[12'hAE2] = 12'hF00;
	mem[12'hAE3] = 12'hF00;
	mem[12'hAE4] = 12'hF00;
	mem[12'hAE5] = 12'hF00;
	mem[12'hAE6] = 12'hF00;
	mem[12'hAE7] = 12'hF00;
	mem[12'hAE8] = 12'hF00;
	mem[12'hAE9] = 12'hF00;
	mem[12'hAEA] = 12'hF00;
	mem[12'hAEB] = 12'hF00;
	mem[12'hAEC] = 12'hF00;
	mem[12'hAED] = 12'hF00;
	mem[12'hAEE] = 12'hF00;
	mem[12'hAEF] = 12'hF00;
	mem[12'hAF0] = 12'hF00;
	mem[12'hAF1] = 12'hF00;
	mem[12'hAF2] = 12'hF00;
	mem[12'hAF3] = 12'hF00;
	mem[12'hAF4] = 12'hF00;
	mem[12'hAF5] = 12'hF00;
	mem[12'hAF6] = 12'hF00;
	mem[12'hAF7] = 12'hF00;
	mem[12'hAF8] = 12'hE22;
	mem[12'hAF9] = 12'hFFF;
	mem[12'hAFA] = 12'hFFF;
	mem[12'hAFB] = 12'hFFF;
	mem[12'hAFC] = 12'hFFF;
	mem[12'hAFD] = 12'hFFF;
	mem[12'hAFE] = 12'hFFF;
	mem[12'hAFF] = 12'hFFF;
	mem[12'hB00] = 12'hFFF;
	mem[12'hB01] = 12'hFFF;
	mem[12'hB02] = 12'hFFF;
	mem[12'hB03] = 12'hFFF;
	mem[12'hB04] = 12'hFFF;
	mem[12'hB05] = 12'hFFF;
	mem[12'hB06] = 12'hFFF;
	mem[12'hB07] = 12'hE22;
	mem[12'hB08] = 12'hF00;
	mem[12'hB09] = 12'hF00;
	mem[12'hB0A] = 12'hF00;
	mem[12'hB0B] = 12'hF00;
	mem[12'hB0C] = 12'hF00;
	mem[12'hB0D] = 12'hF00;
	mem[12'hB0E] = 12'hF00;
	mem[12'hB0F] = 12'hF00;
	mem[12'hB10] = 12'hF00;
	mem[12'hB11] = 12'hF00;
	mem[12'hB12] = 12'hF00;
	mem[12'hB13] = 12'hF00;
	mem[12'hB14] = 12'hF00;
	mem[12'hB15] = 12'hF00;
	mem[12'hB16] = 12'hF00;
	mem[12'hB17] = 12'hF00;
	mem[12'hB18] = 12'hF00;
	mem[12'hB19] = 12'hF00;
	mem[12'hB1A] = 12'hF00;
	mem[12'hB1B] = 12'hF00;
	mem[12'hB1C] = 12'hF00;
	mem[12'hB1D] = 12'hF00;
	mem[12'hB1E] = 12'hF00;
	mem[12'hB1F] = 12'hF00;
	mem[12'hB20] = 12'hF00;
	mem[12'hB21] = 12'hF00;
	mem[12'hB22] = 12'hF00;
	mem[12'hB23] = 12'hF00;
	mem[12'hB24] = 12'hF00;
	mem[12'hB25] = 12'hF00;
	mem[12'hB26] = 12'hF00;
	mem[12'hB27] = 12'hF00;
	mem[12'hB28] = 12'hF00;
	mem[12'hB29] = 12'hF00;
	mem[12'hB2A] = 12'hF00;
	mem[12'hB2B] = 12'hF00;
	mem[12'hB2C] = 12'hF00;
	mem[12'hB2D] = 12'hF00;
	mem[12'hB2E] = 12'hF00;
	mem[12'hB2F] = 12'hF00;
	mem[12'hB30] = 12'hF00;
	mem[12'hB31] = 12'hF00;
	mem[12'hB32] = 12'hF00;
	mem[12'hB33] = 12'hF00;
	mem[12'hB34] = 12'hF00;
	mem[12'hB35] = 12'hF00;
	mem[12'hB36] = 12'hF00;
	mem[12'hB37] = 12'hF00;
	mem[12'hB38] = 12'hE22;
	mem[12'hB39] = 12'hFFF;
	mem[12'hB3A] = 12'hFFF;
	mem[12'hB3B] = 12'hFFF;
	mem[12'hB3C] = 12'hFFF;
	mem[12'hB3D] = 12'hFFF;
	mem[12'hB3E] = 12'hFFF;
	mem[12'hB3F] = 12'hFFF;
	mem[12'hB40] = 12'hFFF;
	mem[12'hB41] = 12'hFFF;
	mem[12'hB42] = 12'hFFF;
	mem[12'hB43] = 12'hFFF;
	mem[12'hB44] = 12'hFFF;
	mem[12'hB45] = 12'hFFF;
	mem[12'hB46] = 12'hFFF;
	mem[12'hB47] = 12'hE22;
	mem[12'hB48] = 12'hF00;
	mem[12'hB49] = 12'hF00;
	mem[12'hB4A] = 12'hF00;
	mem[12'hB4B] = 12'hF00;
	mem[12'hB4C] = 12'hF00;
	mem[12'hB4D] = 12'hF00;
	mem[12'hB4E] = 12'hF00;
	mem[12'hB4F] = 12'hF00;
	mem[12'hB50] = 12'hF00;
	mem[12'hB51] = 12'hF00;
	mem[12'hB52] = 12'hF00;
	mem[12'hB53] = 12'hF00;
	mem[12'hB54] = 12'hF00;
	mem[12'hB55] = 12'hF00;
	mem[12'hB56] = 12'hF00;
	mem[12'hB57] = 12'hF00;
	mem[12'hB58] = 12'hF00;
	mem[12'hB59] = 12'hF00;
	mem[12'hB5A] = 12'hF00;
	mem[12'hB5B] = 12'hF00;
	mem[12'hB5C] = 12'hF00;
	mem[12'hB5D] = 12'hF00;
	mem[12'hB5E] = 12'hF00;
	mem[12'hB5F] = 12'hF00;
	mem[12'hB60] = 12'hF00;
	mem[12'hB61] = 12'hF00;
	mem[12'hB62] = 12'hF00;
	mem[12'hB63] = 12'hF00;
	mem[12'hB64] = 12'hF00;
	mem[12'hB65] = 12'hF00;
	mem[12'hB66] = 12'hF00;
	mem[12'hB67] = 12'hF00;
	mem[12'hB68] = 12'hF00;
	mem[12'hB69] = 12'hF00;
	mem[12'hB6A] = 12'hF00;
	mem[12'hB6B] = 12'hF00;
	mem[12'hB6C] = 12'hF00;
	mem[12'hB6D] = 12'hF00;
	mem[12'hB6E] = 12'hF00;
	mem[12'hB6F] = 12'hF00;
	mem[12'hB70] = 12'hF00;
	mem[12'hB71] = 12'hF00;
	mem[12'hB72] = 12'hF00;
	mem[12'hB73] = 12'hF00;
	mem[12'hB74] = 12'hF00;
	mem[12'hB75] = 12'hF00;
	mem[12'hB76] = 12'hF00;
	mem[12'hB77] = 12'hF00;
	mem[12'hB78] = 12'hE22;
	mem[12'hB79] = 12'hFFF;
	mem[12'hB7A] = 12'hFFF;
	mem[12'hB7B] = 12'hFFF;
	mem[12'hB7C] = 12'hFFF;
	mem[12'hB7D] = 12'hFFF;
	mem[12'hB7E] = 12'hFFF;
	mem[12'hB7F] = 12'hFFF;
	mem[12'hB80] = 12'hFFF;
	mem[12'hB81] = 12'hFFF;
	mem[12'hB82] = 12'hFFF;
	mem[12'hB83] = 12'hFFF;
	mem[12'hB84] = 12'hFFF;
	mem[12'hB85] = 12'hFFF;
	mem[12'hB86] = 12'hFFF;
	mem[12'hB87] = 12'hE22;
	mem[12'hB88] = 12'hF00;
	mem[12'hB89] = 12'hF00;
	mem[12'hB8A] = 12'hF00;
	mem[12'hB8B] = 12'hF00;
	mem[12'hB8C] = 12'hF00;
	mem[12'hB8D] = 12'hF00;
	mem[12'hB8E] = 12'hF00;
	mem[12'hB8F] = 12'hF00;
	mem[12'hB90] = 12'hF00;
	mem[12'hB91] = 12'hF00;
	mem[12'hB92] = 12'hF00;
	mem[12'hB93] = 12'hF00;
	mem[12'hB94] = 12'hF00;
	mem[12'hB95] = 12'hF00;
	mem[12'hB96] = 12'hF00;
	mem[12'hB97] = 12'hF00;
	mem[12'hB98] = 12'hF00;
	mem[12'hB99] = 12'hF00;
	mem[12'hB9A] = 12'hF00;
	mem[12'hB9B] = 12'hF00;
	mem[12'hB9C] = 12'hF00;
	mem[12'hB9D] = 12'hF00;
	mem[12'hB9E] = 12'hF00;
	mem[12'hB9F] = 12'hF00;
	mem[12'hBA0] = 12'hF00;
	mem[12'hBA1] = 12'hF00;
	mem[12'hBA2] = 12'hF00;
	mem[12'hBA3] = 12'hF00;
	mem[12'hBA4] = 12'hF00;
	mem[12'hBA5] = 12'hF00;
	mem[12'hBA6] = 12'hF00;
	mem[12'hBA7] = 12'hF00;
	mem[12'hBA8] = 12'hF00;
	mem[12'hBA9] = 12'hF00;
	mem[12'hBAA] = 12'hF00;
	mem[12'hBAB] = 12'hF00;
	mem[12'hBAC] = 12'hF00;
	mem[12'hBAD] = 12'hF00;
	mem[12'hBAE] = 12'hF00;
	mem[12'hBAF] = 12'hF00;
	mem[12'hBB0] = 12'hF00;
	mem[12'hBB1] = 12'hF00;
	mem[12'hBB2] = 12'hF00;
	mem[12'hBB3] = 12'hF00;
	mem[12'hBB4] = 12'hF00;
	mem[12'hBB5] = 12'hF00;
	mem[12'hBB6] = 12'hF00;
	mem[12'hBB7] = 12'hF00;
	mem[12'hBB8] = 12'hE22;
	mem[12'hBB9] = 12'hFFF;
	mem[12'hBBA] = 12'hFFF;
	mem[12'hBBB] = 12'hFFF;
	mem[12'hBBC] = 12'hFFF;
	mem[12'hBBD] = 12'hFFF;
	mem[12'hBBE] = 12'hFFF;
	mem[12'hBBF] = 12'hFFF;
	mem[12'hBC0] = 12'hFFF;
	mem[12'hBC1] = 12'hFFF;
	mem[12'hBC2] = 12'hFFF;
	mem[12'hBC3] = 12'hFFF;
	mem[12'hBC4] = 12'hFFF;
	mem[12'hBC5] = 12'hFFF;
	mem[12'hBC6] = 12'hFFF;
	mem[12'hBC7] = 12'hE22;
	mem[12'hBC8] = 12'hF00;
	mem[12'hBC9] = 12'hF00;
	mem[12'hBCA] = 12'hF00;
	mem[12'hBCB] = 12'hF00;
	mem[12'hBCC] = 12'hF00;
	mem[12'hBCD] = 12'hF00;
	mem[12'hBCE] = 12'hF00;
	mem[12'hBCF] = 12'hF00;
	mem[12'hBD0] = 12'hF00;
	mem[12'hBD1] = 12'hF00;
	mem[12'hBD2] = 12'hF00;
	mem[12'hBD3] = 12'hF00;
	mem[12'hBD4] = 12'hF00;
	mem[12'hBD5] = 12'hF00;
	mem[12'hBD6] = 12'hF00;
	mem[12'hBD7] = 12'hF00;
	mem[12'hBD8] = 12'hF00;
	mem[12'hBD9] = 12'hF00;
	mem[12'hBDA] = 12'hF00;
	mem[12'hBDB] = 12'hF00;
	mem[12'hBDC] = 12'hF00;
	mem[12'hBDD] = 12'hF00;
	mem[12'hBDE] = 12'hF00;
	mem[12'hBDF] = 12'hF00;
	mem[12'hBE0] = 12'hF00;
	mem[12'hBE1] = 12'hF00;
	mem[12'hBE2] = 12'hF00;
	mem[12'hBE3] = 12'hF00;
	mem[12'hBE4] = 12'hF00;
	mem[12'hBE5] = 12'hF00;
	mem[12'hBE6] = 12'hF00;
	mem[12'hBE7] = 12'hF00;
	mem[12'hBE8] = 12'hF00;
	mem[12'hBE9] = 12'hF00;
	mem[12'hBEA] = 12'hF00;
	mem[12'hBEB] = 12'hF00;
	mem[12'hBEC] = 12'hF00;
	mem[12'hBED] = 12'hF00;
	mem[12'hBEE] = 12'hF00;
	mem[12'hBEF] = 12'hF00;
	mem[12'hBF0] = 12'hF00;
	mem[12'hBF1] = 12'hF00;
	mem[12'hBF2] = 12'hF00;
	mem[12'hBF3] = 12'hF00;
	mem[12'hBF4] = 12'hF00;
	mem[12'hBF5] = 12'hF00;
	mem[12'hBF6] = 12'hF00;
	mem[12'hBF7] = 12'hF00;
	mem[12'hBF8] = 12'hE22;
	mem[12'hBF9] = 12'hFFF;
	mem[12'hBFA] = 12'hFFF;
	mem[12'hBFB] = 12'hFFF;
	mem[12'hBFC] = 12'hFFF;
	mem[12'hBFD] = 12'hFFF;
	mem[12'hBFE] = 12'hFFF;
	mem[12'hBFF] = 12'hFFF;
	mem[12'hC00] = 12'hFFF;
	mem[12'hC01] = 12'hFFF;
	mem[12'hC02] = 12'hFFF;
	mem[12'hC03] = 12'hFFF;
	mem[12'hC04] = 12'hFFF;
	mem[12'hC05] = 12'hFFF;
	mem[12'hC06] = 12'hFFF;
	mem[12'hC07] = 12'hE22;
	mem[12'hC08] = 12'hF00;
	mem[12'hC09] = 12'hF00;
	mem[12'hC0A] = 12'hF00;
	mem[12'hC0B] = 12'hF00;
	mem[12'hC0C] = 12'hF00;
	mem[12'hC0D] = 12'hF00;
	mem[12'hC0E] = 12'hF00;
	mem[12'hC0F] = 12'hF00;
	mem[12'hC10] = 12'hF00;
	mem[12'hC11] = 12'hF00;
	mem[12'hC12] = 12'hF00;
	mem[12'hC13] = 12'hF00;
	mem[12'hC14] = 12'hF00;
	mem[12'hC15] = 12'hF00;
	mem[12'hC16] = 12'hF00;
	mem[12'hC17] = 12'hF00;
	mem[12'hC18] = 12'hF00;
	mem[12'hC19] = 12'hF00;
	mem[12'hC1A] = 12'hF00;
	mem[12'hC1B] = 12'hF00;
	mem[12'hC1C] = 12'hF00;
	mem[12'hC1D] = 12'hF00;
	mem[12'hC1E] = 12'hF00;
	mem[12'hC1F] = 12'hF00;
	mem[12'hC20] = 12'hF00;
	mem[12'hC21] = 12'hF00;
	mem[12'hC22] = 12'hF00;
	mem[12'hC23] = 12'hF00;
	mem[12'hC24] = 12'hF00;
	mem[12'hC25] = 12'hF00;
	mem[12'hC26] = 12'hF00;
	mem[12'hC27] = 12'hF00;
	mem[12'hC28] = 12'hF00;
	mem[12'hC29] = 12'hF00;
	mem[12'hC2A] = 12'hF00;
	mem[12'hC2B] = 12'hF00;
	mem[12'hC2C] = 12'hF00;
	mem[12'hC2D] = 12'hF00;
	mem[12'hC2E] = 12'hF00;
	mem[12'hC2F] = 12'hF00;
	mem[12'hC30] = 12'hF00;
	mem[12'hC31] = 12'hF00;
	mem[12'hC32] = 12'hF00;
	mem[12'hC33] = 12'hF00;
	mem[12'hC34] = 12'hF00;
	mem[12'hC35] = 12'hF00;
	mem[12'hC36] = 12'hF00;
	mem[12'hC37] = 12'hF00;
	mem[12'hC38] = 12'hE22;
	mem[12'hC39] = 12'hFFF;
	mem[12'hC3A] = 12'hFFF;
	mem[12'hC3B] = 12'hFFF;
	mem[12'hC3C] = 12'hFFF;
	mem[12'hC3D] = 12'hFFF;
	mem[12'hC3E] = 12'hFFF;
	mem[12'hC3F] = 12'hFFF;
	mem[12'hC40] = 12'hFFF;
	mem[12'hC41] = 12'hFFF;
	mem[12'hC42] = 12'hFFF;
	mem[12'hC43] = 12'hFFF;
	mem[12'hC44] = 12'hFFF;
	mem[12'hC45] = 12'hFFF;
	mem[12'hC46] = 12'hFFF;
	mem[12'hC47] = 12'hE22;
	mem[12'hC48] = 12'hF00;
	mem[12'hC49] = 12'hF00;
	mem[12'hC4A] = 12'hF00;
	mem[12'hC4B] = 12'hF00;
	mem[12'hC4C] = 12'hF00;
	mem[12'hC4D] = 12'hF00;
	mem[12'hC4E] = 12'hF00;
	mem[12'hC4F] = 12'hF00;
	mem[12'hC50] = 12'hF00;
	mem[12'hC51] = 12'hF00;
	mem[12'hC52] = 12'hF00;
	mem[12'hC53] = 12'hF00;
	mem[12'hC54] = 12'hF00;
	mem[12'hC55] = 12'hF00;
	mem[12'hC56] = 12'hF00;
	mem[12'hC57] = 12'hF00;
	mem[12'hC58] = 12'hF00;
	mem[12'hC59] = 12'hF00;
	mem[12'hC5A] = 12'hF00;
	mem[12'hC5B] = 12'hF00;
	mem[12'hC5C] = 12'hF00;
	mem[12'hC5D] = 12'hF00;
	mem[12'hC5E] = 12'hF00;
	mem[12'hC5F] = 12'hF00;
	mem[12'hC60] = 12'hF00;
	mem[12'hC61] = 12'hF00;
	mem[12'hC62] = 12'hF00;
	mem[12'hC63] = 12'hF00;
	mem[12'hC64] = 12'hF00;
	mem[12'hC65] = 12'hF00;
	mem[12'hC66] = 12'hF00;
	mem[12'hC67] = 12'hF00;
	mem[12'hC68] = 12'hF00;
	mem[12'hC69] = 12'hF00;
	mem[12'hC6A] = 12'hF00;
	mem[12'hC6B] = 12'hF00;
	mem[12'hC6C] = 12'hF00;
	mem[12'hC6D] = 12'hF00;
	mem[12'hC6E] = 12'hF00;
	mem[12'hC6F] = 12'hF00;
	mem[12'hC70] = 12'hF00;
	mem[12'hC71] = 12'hF00;
	mem[12'hC72] = 12'hF00;
	mem[12'hC73] = 12'hF00;
	mem[12'hC74] = 12'hF00;
	mem[12'hC75] = 12'hF00;
	mem[12'hC76] = 12'hF00;
	mem[12'hC77] = 12'hF00;
	mem[12'hC78] = 12'hE22;
	mem[12'hC79] = 12'hFFF;
	mem[12'hC7A] = 12'hFFF;
	mem[12'hC7B] = 12'hFFF;
	mem[12'hC7C] = 12'hFFF;
	mem[12'hC7D] = 12'hFFF;
	mem[12'hC7E] = 12'hFFF;
	mem[12'hC7F] = 12'hFFF;
	mem[12'hC80] = 12'hFFF;
	mem[12'hC81] = 12'hFFF;
	mem[12'hC82] = 12'hFFF;
	mem[12'hC83] = 12'hFFF;
	mem[12'hC84] = 12'hFFF;
	mem[12'hC85] = 12'hFFF;
	mem[12'hC86] = 12'hFFF;
	mem[12'hC87] = 12'hE22;
	mem[12'hC88] = 12'hF00;
	mem[12'hC89] = 12'hF00;
	mem[12'hC8A] = 12'hF00;
	mem[12'hC8B] = 12'hF00;
	mem[12'hC8C] = 12'hF00;
	mem[12'hC8D] = 12'hF00;
	mem[12'hC8E] = 12'hF00;
	mem[12'hC8F] = 12'hF00;
	mem[12'hC90] = 12'hF00;
	mem[12'hC91] = 12'hF00;
	mem[12'hC92] = 12'hF00;
	mem[12'hC93] = 12'hF00;
	mem[12'hC94] = 12'hF00;
	mem[12'hC95] = 12'hF00;
	mem[12'hC96] = 12'hF00;
	mem[12'hC97] = 12'hF00;
	mem[12'hC98] = 12'hF00;
	mem[12'hC99] = 12'hF00;
	mem[12'hC9A] = 12'hF00;
	mem[12'hC9B] = 12'hF00;
	mem[12'hC9C] = 12'hF00;
	mem[12'hC9D] = 12'hF00;
	mem[12'hC9E] = 12'hF00;
	mem[12'hC9F] = 12'hF00;
	mem[12'hCA0] = 12'hF00;
	mem[12'hCA1] = 12'hF00;
	mem[12'hCA2] = 12'hF00;
	mem[12'hCA3] = 12'hF00;
	mem[12'hCA4] = 12'hF00;
	mem[12'hCA5] = 12'hF00;
	mem[12'hCA6] = 12'hF00;
	mem[12'hCA7] = 12'hF00;
	mem[12'hCA8] = 12'hF00;
	mem[12'hCA9] = 12'hF00;
	mem[12'hCAA] = 12'hF00;
	mem[12'hCAB] = 12'hF00;
	mem[12'hCAC] = 12'hF00;
	mem[12'hCAD] = 12'hF00;
	mem[12'hCAE] = 12'hF00;
	mem[12'hCAF] = 12'hF00;
	mem[12'hCB0] = 12'hF00;
	mem[12'hCB1] = 12'hF00;
	mem[12'hCB2] = 12'hF00;
	mem[12'hCB3] = 12'hF00;
	mem[12'hCB4] = 12'hF00;
	mem[12'hCB5] = 12'hF00;
	mem[12'hCB6] = 12'hF00;
	mem[12'hCB7] = 12'hF00;
	mem[12'hCB8] = 12'hE22;
	mem[12'hCB9] = 12'hFFF;
	mem[12'hCBA] = 12'hFFF;
	mem[12'hCBB] = 12'hFFF;
	mem[12'hCBC] = 12'hFFF;
	mem[12'hCBD] = 12'hFFF;
	mem[12'hCBE] = 12'hFFF;
	mem[12'hCBF] = 12'hFFF;
	mem[12'hCC0] = 12'hFFF;
	mem[12'hCC1] = 12'hFFF;
	mem[12'hCC2] = 12'hFFF;
	mem[12'hCC3] = 12'hFFF;
	mem[12'hCC4] = 12'hFFF;
	mem[12'hCC5] = 12'hFFF;
	mem[12'hCC6] = 12'hFFF;
	mem[12'hCC7] = 12'hE22;
	mem[12'hCC8] = 12'hF00;
	mem[12'hCC9] = 12'hF00;
	mem[12'hCCA] = 12'hF00;
	mem[12'hCCB] = 12'hF00;
	mem[12'hCCC] = 12'hF00;
	mem[12'hCCD] = 12'hF00;
	mem[12'hCCE] = 12'hF00;
	mem[12'hCCF] = 12'hF00;
	mem[12'hCD0] = 12'hF00;
	mem[12'hCD1] = 12'hF00;
	mem[12'hCD2] = 12'hF00;
	mem[12'hCD3] = 12'hF00;
	mem[12'hCD4] = 12'hF00;
	mem[12'hCD5] = 12'hF00;
	mem[12'hCD6] = 12'hF00;
	mem[12'hCD7] = 12'hF00;
	mem[12'hCD8] = 12'hF00;
	mem[12'hCD9] = 12'hF00;
	mem[12'hCDA] = 12'hF00;
	mem[12'hCDB] = 12'hF00;
	mem[12'hCDC] = 12'hF00;
	mem[12'hCDD] = 12'hF00;
	mem[12'hCDE] = 12'hF00;
	mem[12'hCDF] = 12'hF00;
	mem[12'hCE0] = 12'hF00;
	mem[12'hCE1] = 12'hF00;
	mem[12'hCE2] = 12'hF00;
	mem[12'hCE3] = 12'hF00;
	mem[12'hCE4] = 12'hF00;
	mem[12'hCE5] = 12'hF00;
	mem[12'hCE6] = 12'hF00;
	mem[12'hCE7] = 12'hF00;
	mem[12'hCE8] = 12'hF00;
	mem[12'hCE9] = 12'hF00;
	mem[12'hCEA] = 12'hF00;
	mem[12'hCEB] = 12'hF00;
	mem[12'hCEC] = 12'hF00;
	mem[12'hCED] = 12'hF00;
	mem[12'hCEE] = 12'hF00;
	mem[12'hCEF] = 12'hF00;
	mem[12'hCF0] = 12'hF00;
	mem[12'hCF1] = 12'hF00;
	mem[12'hCF2] = 12'hF00;
	mem[12'hCF3] = 12'hF00;
	mem[12'hCF4] = 12'hF00;
	mem[12'hCF5] = 12'hF00;
	mem[12'hCF6] = 12'hF00;
	mem[12'hCF7] = 12'hF00;
	mem[12'hCF8] = 12'hE22;
	mem[12'hCF9] = 12'hFFF;
	mem[12'hCFA] = 12'hFFF;
	mem[12'hCFB] = 12'hFFF;
	mem[12'hCFC] = 12'hFFF;
	mem[12'hCFD] = 12'hFFF;
	mem[12'hCFE] = 12'hFFF;
	mem[12'hCFF] = 12'hFFF;
	mem[12'hD00] = 12'hFFF;
	mem[12'hD01] = 12'hFFF;
	mem[12'hD02] = 12'hFFF;
	mem[12'hD03] = 12'hFFF;
	mem[12'hD04] = 12'hFFF;
	mem[12'hD05] = 12'hFFF;
	mem[12'hD06] = 12'hFFF;
	mem[12'hD07] = 12'hE22;
	mem[12'hD08] = 12'hF00;
	mem[12'hD09] = 12'hF00;
	mem[12'hD0A] = 12'hF00;
	mem[12'hD0B] = 12'hF00;
	mem[12'hD0C] = 12'hF00;
	mem[12'hD0D] = 12'hF00;
	mem[12'hD0E] = 12'hF00;
	mem[12'hD0F] = 12'hF00;
	mem[12'hD10] = 12'hF00;
	mem[12'hD11] = 12'hF00;
	mem[12'hD12] = 12'hF00;
	mem[12'hD13] = 12'hF00;
	mem[12'hD14] = 12'hF00;
	mem[12'hD15] = 12'hF00;
	mem[12'hD16] = 12'hF00;
	mem[12'hD17] = 12'hF00;
	mem[12'hD18] = 12'hF00;
	mem[12'hD19] = 12'hF00;
	mem[12'hD1A] = 12'hF00;
	mem[12'hD1B] = 12'hF00;
	mem[12'hD1C] = 12'hF00;
	mem[12'hD1D] = 12'hF00;
	mem[12'hD1E] = 12'hF00;
	mem[12'hD1F] = 12'hF00;
	mem[12'hD20] = 12'hF00;
	mem[12'hD21] = 12'hF00;
	mem[12'hD22] = 12'hF00;
	mem[12'hD23] = 12'hF00;
	mem[12'hD24] = 12'hF00;
	mem[12'hD25] = 12'hF00;
	mem[12'hD26] = 12'hF00;
	mem[12'hD27] = 12'hF00;
	mem[12'hD28] = 12'hF00;
	mem[12'hD29] = 12'hF00;
	mem[12'hD2A] = 12'hF00;
	mem[12'hD2B] = 12'hF00;
	mem[12'hD2C] = 12'hF00;
	mem[12'hD2D] = 12'hF00;
	mem[12'hD2E] = 12'hF00;
	mem[12'hD2F] = 12'hF00;
	mem[12'hD30] = 12'hF00;
	mem[12'hD31] = 12'hF00;
	mem[12'hD32] = 12'hF00;
	mem[12'hD33] = 12'hF00;
	mem[12'hD34] = 12'hF00;
	mem[12'hD35] = 12'hF00;
	mem[12'hD36] = 12'hF00;
	mem[12'hD37] = 12'hF00;
	mem[12'hD38] = 12'hE22;
	mem[12'hD39] = 12'hFFF;
	mem[12'hD3A] = 12'hFFF;
	mem[12'hD3B] = 12'hFFF;
	mem[12'hD3C] = 12'hFFF;
	mem[12'hD3D] = 12'hFFF;
	mem[12'hD3E] = 12'hFFF;
	mem[12'hD3F] = 12'hFFF;
	mem[12'hD40] = 12'hFFF;
	mem[12'hD41] = 12'hFFF;
	mem[12'hD42] = 12'hFFF;
	mem[12'hD43] = 12'hFFF;
	mem[12'hD44] = 12'hFFF;
	mem[12'hD45] = 12'hFFF;
	mem[12'hD46] = 12'hFFF;
	mem[12'hD47] = 12'hE22;
	mem[12'hD48] = 12'hF00;
	mem[12'hD49] = 12'hF00;
	mem[12'hD4A] = 12'hF00;
	mem[12'hD4B] = 12'hF00;
	mem[12'hD4C] = 12'hF00;
	mem[12'hD4D] = 12'hF00;
	mem[12'hD4E] = 12'hF00;
	mem[12'hD4F] = 12'hF00;
	mem[12'hD50] = 12'hE22;
	mem[12'hD51] = 12'hE22;
	mem[12'hD52] = 12'hE22;
	mem[12'hD53] = 12'hF00;
	mem[12'hD54] = 12'hF00;
	mem[12'hD55] = 12'hF00;
	mem[12'hD56] = 12'hF00;
	mem[12'hD57] = 12'hF00;
	mem[12'hD58] = 12'hF00;
	mem[12'hD59] = 12'hF00;
	mem[12'hD5A] = 12'hF00;
	mem[12'hD5B] = 12'hF00;
	mem[12'hD5C] = 12'hF00;
	mem[12'hD5D] = 12'hF00;
	mem[12'hD5E] = 12'hE22;
	mem[12'hD5F] = 12'hE22;
	mem[12'hD60] = 12'hE22;
	mem[12'hD61] = 12'hE22;
	mem[12'hD62] = 12'hF00;
	mem[12'hD63] = 12'hF00;
	mem[12'hD64] = 12'hF00;
	mem[12'hD65] = 12'hF00;
	mem[12'hD66] = 12'hF00;
	mem[12'hD67] = 12'hF00;
	mem[12'hD68] = 12'hF00;
	mem[12'hD69] = 12'hF00;
	mem[12'hD6A] = 12'hF00;
	mem[12'hD6B] = 12'hF00;
	mem[12'hD6C] = 12'hF00;
	mem[12'hD6D] = 12'hF00;
	mem[12'hD6E] = 12'hE22;
	mem[12'hD6F] = 12'hE22;
	mem[12'hD70] = 12'hE22;
	mem[12'hD71] = 12'hF00;
	mem[12'hD72] = 12'hF00;
	mem[12'hD73] = 12'hF00;
	mem[12'hD74] = 12'hF00;
	mem[12'hD75] = 12'hF00;
	mem[12'hD76] = 12'hF00;
	mem[12'hD77] = 12'hF00;
	mem[12'hD78] = 12'hE22;
	mem[12'hD79] = 12'hFFF;
	mem[12'hD7A] = 12'hFFF;
	mem[12'hD7B] = 12'hFFF;
	mem[12'hD7C] = 12'hFFF;
	mem[12'hD7D] = 12'hFFF;
	mem[12'hD7E] = 12'hFFF;
	mem[12'hD7F] = 12'hFFF;
	mem[12'hD80] = 12'hFFF;
	mem[12'hD81] = 12'hFFF;
	mem[12'hD82] = 12'hFFF;
	mem[12'hD83] = 12'hFFF;
	mem[12'hD84] = 12'hFFF;
	mem[12'hD85] = 12'hFFF;
	mem[12'hD86] = 12'hFFF;
	mem[12'hD87] = 12'hF00;
	mem[12'hD88] = 12'hF00;
	mem[12'hD89] = 12'hF00;
	mem[12'hD8A] = 12'hF00;
	mem[12'hD8B] = 12'hF00;
	mem[12'hD8C] = 12'hF00;
	mem[12'hD8D] = 12'hF00;
	mem[12'hD8E] = 12'hF00;
	mem[12'hD8F] = 12'hF00;
	mem[12'hD90] = 12'hFFF;
	mem[12'hD91] = 12'hFFF;
	mem[12'hD92] = 12'hFFF;
	mem[12'hD93] = 12'hE22;
	mem[12'hD94] = 12'hF00;
	mem[12'hD95] = 12'hF00;
	mem[12'hD96] = 12'hF00;
	mem[12'hD97] = 12'hF00;
	mem[12'hD98] = 12'hF00;
	mem[12'hD99] = 12'hF00;
	mem[12'hD9A] = 12'hF00;
	mem[12'hD9B] = 12'hF00;
	mem[12'hD9C] = 12'hF00;
	mem[12'hD9D] = 12'hE22;
	mem[12'hD9E] = 12'hFFF;
	mem[12'hD9F] = 12'hFFF;
	mem[12'hDA0] = 12'hFFF;
	mem[12'hDA1] = 12'hFFF;
	mem[12'hDA2] = 12'hE22;
	mem[12'hDA3] = 12'hF00;
	mem[12'hDA4] = 12'hF00;
	mem[12'hDA5] = 12'hF00;
	mem[12'hDA6] = 12'hF00;
	mem[12'hDA7] = 12'hF00;
	mem[12'hDA8] = 12'hF00;
	mem[12'hDA9] = 12'hF00;
	mem[12'hDAA] = 12'hF00;
	mem[12'hDAB] = 12'hF00;
	mem[12'hDAC] = 12'hF00;
	mem[12'hDAD] = 12'hE22;
	mem[12'hDAE] = 12'hFFF;
	mem[12'hDAF] = 12'hFFF;
	mem[12'hDB0] = 12'hFFF;
	mem[12'hDB1] = 12'hF00;
	mem[12'hDB2] = 12'hF00;
	mem[12'hDB3] = 12'hF00;
	mem[12'hDB4] = 12'hF00;
	mem[12'hDB5] = 12'hF00;
	mem[12'hDB6] = 12'hF00;
	mem[12'hDB7] = 12'hF00;
	mem[12'hDB8] = 12'hE22;
	mem[12'hDB9] = 12'hFFF;
	mem[12'hDBA] = 12'hFFF;
	mem[12'hDBB] = 12'hFFF;
	mem[12'hDBC] = 12'hFFF;
	mem[12'hDBD] = 12'hFFF;
	mem[12'hDBE] = 12'hFFF;
	mem[12'hDBF] = 12'hFFF;
	mem[12'hDC0] = 12'hFFF;
	mem[12'hDC1] = 12'hFFF;
	mem[12'hDC2] = 12'hFFF;
	mem[12'hDC3] = 12'hFFF;
	mem[12'hDC4] = 12'hFFF;
	mem[12'hDC5] = 12'hFFF;
	mem[12'hDC6] = 12'hFFF;
	mem[12'hDC7] = 12'hF00;
	mem[12'hDC8] = 12'hF00;
	mem[12'hDC9] = 12'hF00;
	mem[12'hDCA] = 12'hF00;
	mem[12'hDCB] = 12'hF00;
	mem[12'hDCC] = 12'hF00;
	mem[12'hDCD] = 12'hE22;
	mem[12'hDCE] = 12'hF00;
	mem[12'hDCF] = 12'hFFF;
	mem[12'hDD0] = 12'hFFF;
	mem[12'hDD1] = 12'hFFF;
	mem[12'hDD2] = 12'hFFF;
	mem[12'hDD3] = 12'hFFF;
	mem[12'hDD4] = 12'hE22;
	mem[12'hDD5] = 12'hF00;
	mem[12'hDD6] = 12'hF00;
	mem[12'hDD7] = 12'hF00;
	mem[12'hDD8] = 12'hF00;
	mem[12'hDD9] = 12'hF00;
	mem[12'hDDA] = 12'hF00;
	mem[12'hDDB] = 12'hF00;
	mem[12'hDDC] = 12'hE22;
	mem[12'hDDD] = 12'hFFF;
	mem[12'hDDE] = 12'hFFF;
	mem[12'hDDF] = 12'hFFF;
	mem[12'hDE0] = 12'hFFF;
	mem[12'hDE1] = 12'hFFF;
	mem[12'hDE2] = 12'hFFF;
	mem[12'hDE3] = 12'hE22;
	mem[12'hDE4] = 12'hF00;
	mem[12'hDE5] = 12'hF00;
	mem[12'hDE6] = 12'hF00;
	mem[12'hDE7] = 12'hF00;
	mem[12'hDE8] = 12'hF00;
	mem[12'hDE9] = 12'hF00;
	mem[12'hDEA] = 12'hF00;
	mem[12'hDEB] = 12'hF00;
	mem[12'hDEC] = 12'hE22;
	mem[12'hDED] = 12'hFFF;
	mem[12'hDEE] = 12'hFFF;
	mem[12'hDEF] = 12'hFFF;
	mem[12'hDF0] = 12'hFFF;
	mem[12'hDF1] = 12'hFFF;
	mem[12'hDF2] = 12'hF00;
	mem[12'hDF3] = 12'hF00;
	mem[12'hDF4] = 12'hF00;
	mem[12'hDF5] = 12'hF00;
	mem[12'hDF6] = 12'hF00;
	mem[12'hDF7] = 12'hF00;
	mem[12'hDF8] = 12'hF00;
	mem[12'hDF9] = 12'hFFF;
	mem[12'hDFA] = 12'hFFF;
	mem[12'hDFB] = 12'hFFF;
	mem[12'hDFC] = 12'hFFF;
	mem[12'hDFD] = 12'hFFF;
	mem[12'hDFE] = 12'hFFF;
	mem[12'hDFF] = 12'hFFF;
	mem[12'hE00] = 12'hFFF;
	mem[12'hE01] = 12'hFFF;
	mem[12'hE02] = 12'hFFF;
	mem[12'hE03] = 12'hFFF;
	mem[12'hE04] = 12'hFFF;
	mem[12'hE05] = 12'hFFF;
	mem[12'hE06] = 12'hFFF;
	mem[12'hE07] = 12'hF00;
	mem[12'hE08] = 12'hF00;
	mem[12'hE09] = 12'hF00;
	mem[12'hE0A] = 12'hF00;
	mem[12'hE0B] = 12'hF00;
	mem[12'hE0C] = 12'hE22;
	mem[12'hE0D] = 12'hFFF;
	mem[12'hE0E] = 12'hFFF;
	mem[12'hE0F] = 12'hFFF;
	mem[12'hE10] = 12'hFFF;
	mem[12'hE11] = 12'hFFF;
	mem[12'hE12] = 12'hFFF;
	mem[12'hE13] = 12'hFFF;
	mem[12'hE14] = 12'hFFF;
	mem[12'hE15] = 12'hE22;
	mem[12'hE16] = 12'hF00;
	mem[12'hE17] = 12'hF00;
	mem[12'hE18] = 12'hF00;
	mem[12'hE19] = 12'hF00;
	mem[12'hE1A] = 12'hF00;
	mem[12'hE1B] = 12'hE22;
	mem[12'hE1C] = 12'hFFF;
	mem[12'hE1D] = 12'hFFF;
	mem[12'hE1E] = 12'hFFF;
	mem[12'hE1F] = 12'hFFF;
	mem[12'hE20] = 12'hFFF;
	mem[12'hE21] = 12'hFFF;
	mem[12'hE22] = 12'hFFF;
	mem[12'hE23] = 12'hFFF;
	mem[12'hE24] = 12'hE22;
	mem[12'hE25] = 12'hF00;
	mem[12'hE26] = 12'hF00;
	mem[12'hE27] = 12'hF00;
	mem[12'hE28] = 12'hF00;
	mem[12'hE29] = 12'hF00;
	mem[12'hE2A] = 12'hF00;
	mem[12'hE2B] = 12'hE22;
	mem[12'hE2C] = 12'hFFF;
	mem[12'hE2D] = 12'hFFF;
	mem[12'hE2E] = 12'hFFF;
	mem[12'hE2F] = 12'hFFF;
	mem[12'hE30] = 12'hFFF;
	mem[12'hE31] = 12'hFFF;
	mem[12'hE32] = 12'hFFF;
	mem[12'hE33] = 12'hF00;
	mem[12'hE34] = 12'hF00;
	mem[12'hE35] = 12'hF00;
	mem[12'hE36] = 12'hF00;
	mem[12'hE37] = 12'hF00;
	mem[12'hE38] = 12'hF00;
	mem[12'hE39] = 12'hFFF;
	mem[12'hE3A] = 12'hFFF;
	mem[12'hE3B] = 12'hFFF;
	mem[12'hE3C] = 12'hFFF;
	mem[12'hE3D] = 12'hFFF;
	mem[12'hE3E] = 12'hFFF;
	mem[12'hE3F] = 12'hFFF;
	mem[12'hE40] = 12'hFFF;
	mem[12'hE41] = 12'hFFF;
	mem[12'hE42] = 12'hFFF;
	mem[12'hE43] = 12'hFFF;
	mem[12'hE44] = 12'hFFF;
	mem[12'hE45] = 12'hFFF;
	mem[12'hE46] = 12'hFFF;
	mem[12'hE47] = 12'hFFF;
	mem[12'hE48] = 12'hF00;
	mem[12'hE49] = 12'hF00;
	mem[12'hE4A] = 12'hF00;
	mem[12'hE4B] = 12'hE22;
	mem[12'hE4C] = 12'hFFF;
	mem[12'hE4D] = 12'hFFF;
	mem[12'hE4E] = 12'hFFF;
	mem[12'hE4F] = 12'hFFF;
	mem[12'hE50] = 12'hFFF;
	mem[12'hE51] = 12'hFFF;
	mem[12'hE52] = 12'hFFF;
	mem[12'hE53] = 12'hFFF;
	mem[12'hE54] = 12'hFFF;
	mem[12'hE55] = 12'hFFF;
	mem[12'hE56] = 12'hE22;
	mem[12'hE57] = 12'hF00;
	mem[12'hE58] = 12'hF00;
	mem[12'hE59] = 12'hF00;
	mem[12'hE5A] = 12'hF00;
	mem[12'hE5B] = 12'hF00;
	mem[12'hE5C] = 12'hFFF;
	mem[12'hE5D] = 12'hFFF;
	mem[12'hE5E] = 12'hFFF;
	mem[12'hE5F] = 12'hFFF;
	mem[12'hE60] = 12'hFFF;
	mem[12'hE61] = 12'hFFF;
	mem[12'hE62] = 12'hFFF;
	mem[12'hE63] = 12'hFFF;
	mem[12'hE64] = 12'hFFF;
	mem[12'hE65] = 12'hE22;
	mem[12'hE66] = 12'hF00;
	mem[12'hE67] = 12'hF00;
	mem[12'hE68] = 12'hF00;
	mem[12'hE69] = 12'hF00;
	mem[12'hE6A] = 12'hE22;
	mem[12'hE6B] = 12'hFFF;
	mem[12'hE6C] = 12'hFFF;
	mem[12'hE6D] = 12'hFFF;
	mem[12'hE6E] = 12'hFFF;
	mem[12'hE6F] = 12'hFFF;
	mem[12'hE70] = 12'hFFF;
	mem[12'hE71] = 12'hFFF;
	mem[12'hE72] = 12'hFFF;
	mem[12'hE73] = 12'hFFF;
	mem[12'hE74] = 12'hE22;
	mem[12'hE75] = 12'hF00;
	mem[12'hE76] = 12'hF00;
	mem[12'hE77] = 12'hF00;
	mem[12'hE78] = 12'hF00;
	mem[12'hE79] = 12'hFFF;
	mem[12'hE7A] = 12'hFFF;
	mem[12'hE7B] = 12'hFFF;
	mem[12'hE7C] = 12'hFFF;
	mem[12'hE7D] = 12'hFFF;
	mem[12'hE7E] = 12'hFFF;
	mem[12'hE7F] = 12'hFFF;
	mem[12'hE80] = 12'hFFF;
	mem[12'hE81] = 12'hFFF;
	mem[12'hE82] = 12'hFFF;
	mem[12'hE83] = 12'hFFF;
	mem[12'hE84] = 12'hFFF;
	mem[12'hE85] = 12'hFFF;
	mem[12'hE86] = 12'hFFF;
	mem[12'hE87] = 12'hFFF;
	mem[12'hE88] = 12'hE22;
	mem[12'hE89] = 12'hF00;
	mem[12'hE8A] = 12'hE22;
	mem[12'hE8B] = 12'hFFF;
	mem[12'hE8C] = 12'hFFF;
	mem[12'hE8D] = 12'hFFF;
	mem[12'hE8E] = 12'hFFF;
	mem[12'hE8F] = 12'hFFF;
	mem[12'hE90] = 12'hFFF;
	mem[12'hE91] = 12'hFFF;
	mem[12'hE92] = 12'hFFF;
	mem[12'hE93] = 12'hFFF;
	mem[12'hE94] = 12'hFFF;
	mem[12'hE95] = 12'hFFF;
	mem[12'hE96] = 12'hFFF;
	mem[12'hE97] = 12'hE22;
	mem[12'hE98] = 12'hF00;
	mem[12'hE99] = 12'hF00;
	mem[12'hE9A] = 12'hF00;
	mem[12'hE9B] = 12'hFFF;
	mem[12'hE9C] = 12'hFFF;
	mem[12'hE9D] = 12'hFFF;
	mem[12'hE9E] = 12'hFFF;
	mem[12'hE9F] = 12'hFFF;
	mem[12'hEA0] = 12'hFFF;
	mem[12'hEA1] = 12'hFFF;
	mem[12'hEA2] = 12'hFFF;
	mem[12'hEA3] = 12'hFFF;
	mem[12'hEA4] = 12'hFFF;
	mem[12'hEA5] = 12'hFFF;
	mem[12'hEA6] = 12'hE22;
	mem[12'hEA7] = 12'hF00;
	mem[12'hEA8] = 12'hF00;
	mem[12'hEA9] = 12'hE22;
	mem[12'hEAA] = 12'hFFF;
	mem[12'hEAB] = 12'hFFF;
	mem[12'hEAC] = 12'hFFF;
	mem[12'hEAD] = 12'hFFF;
	mem[12'hEAE] = 12'hFFF;
	mem[12'hEAF] = 12'hFFF;
	mem[12'hEB0] = 12'hFFF;
	mem[12'hEB1] = 12'hFFF;
	mem[12'hEB2] = 12'hFFF;
	mem[12'hEB3] = 12'hFFF;
	mem[12'hEB4] = 12'hFFF;
	mem[12'hEB5] = 12'hE22;
	mem[12'hEB6] = 12'hF00;
	mem[12'hEB7] = 12'hE22;
	mem[12'hEB8] = 12'hFFF;
	mem[12'hEB9] = 12'hFFF;
	mem[12'hEBA] = 12'hFFF;
	mem[12'hEBB] = 12'hFFF;
	mem[12'hEBC] = 12'hFFF;
	mem[12'hEBD] = 12'hFFF;
	mem[12'hEBE] = 12'hFFF;
	mem[12'hEBF] = 12'hFFF;
	mem[12'hEC0] = 12'hFFF;
	mem[12'hEC1] = 12'hFFF;
	mem[12'hEC2] = 12'hFFF;
	mem[12'hEC3] = 12'hFFF;
	mem[12'hEC4] = 12'hFFF;
	mem[12'hEC5] = 12'hFFF;
	mem[12'hEC6] = 12'hFFF;
	mem[12'hEC7] = 12'hFFF;
	mem[12'hEC8] = 12'hFFF;
	mem[12'hEC9] = 12'hFFF;
	mem[12'hECA] = 12'hFFF;
	mem[12'hECB] = 12'hFFF;
	mem[12'hECC] = 12'hFFF;
	mem[12'hECD] = 12'hFFF;
	mem[12'hECE] = 12'hFFF;
	mem[12'hECF] = 12'hFFF;
	mem[12'hED0] = 12'hFFF;
	mem[12'hED1] = 12'hFFF;
	mem[12'hED2] = 12'hFFF;
	mem[12'hED3] = 12'hFFF;
	mem[12'hED4] = 12'hFFF;
	mem[12'hED5] = 12'hFFF;
	mem[12'hED6] = 12'hFFF;
	mem[12'hED7] = 12'hFFF;
	mem[12'hED8] = 12'hFFF;
	mem[12'hED9] = 12'hFFF;
	mem[12'hEDA] = 12'hFFF;
	mem[12'hEDB] = 12'hFFF;
	mem[12'hEDC] = 12'hFFF;
	mem[12'hEDD] = 12'hFFF;
	mem[12'hEDE] = 12'hFFF;
	mem[12'hEDF] = 12'hFFF;
	mem[12'hEE0] = 12'hFFF;
	mem[12'hEE1] = 12'hFFF;
	mem[12'hEE2] = 12'hFFF;
	mem[12'hEE3] = 12'hFFF;
	mem[12'hEE4] = 12'hFFF;
	mem[12'hEE5] = 12'hFFF;
	mem[12'hEE6] = 12'hFFF;
	mem[12'hEE7] = 12'hFFF;
	mem[12'hEE8] = 12'hFFF;
	mem[12'hEE9] = 12'hFFF;
	mem[12'hEEA] = 12'hFFF;
	mem[12'hEEB] = 12'hFFF;
	mem[12'hEEC] = 12'hFFF;
	mem[12'hEED] = 12'hFFF;
	mem[12'hEEE] = 12'hFFF;
	mem[12'hEEF] = 12'hFFF;
	mem[12'hEF0] = 12'hFFF;
	mem[12'hEF1] = 12'hFFF;
	mem[12'hEF2] = 12'hFFF;
	mem[12'hEF3] = 12'hFFF;
	mem[12'hEF4] = 12'hFFF;
	mem[12'hEF5] = 12'hFFF;
	mem[12'hEF6] = 12'hFFF;
	mem[12'hEF7] = 12'hFFF;
	mem[12'hEF8] = 12'hFFF;
	mem[12'hEF9] = 12'hFFF;
	mem[12'hEFA] = 12'hFFF;
	mem[12'hEFB] = 12'hFFF;
	mem[12'hEFC] = 12'hFFF;
	mem[12'hEFD] = 12'hFFF;
	mem[12'hEFE] = 12'hFFF;
	mem[12'hEFF] = 12'hFFF;
	mem[12'hF00] = 12'hFFF;
	mem[12'hF01] = 12'hFFF;
	mem[12'hF02] = 12'hFFF;
	mem[12'hF03] = 12'hFFF;
	mem[12'hF04] = 12'hFFF;
	mem[12'hF05] = 12'hFFF;
	mem[12'hF06] = 12'hFFF;
	mem[12'hF07] = 12'hFFF;
	mem[12'hF08] = 12'hFFF;
	mem[12'hF09] = 12'hFFF;
	mem[12'hF0A] = 12'hFFF;
	mem[12'hF0B] = 12'hFFF;
	mem[12'hF0C] = 12'hFFF;
	mem[12'hF0D] = 12'hFFF;
	mem[12'hF0E] = 12'hFFF;
	mem[12'hF0F] = 12'hFFF;
	mem[12'hF10] = 12'hFFF;
	mem[12'hF11] = 12'hFFF;
	mem[12'hF12] = 12'hFFF;
	mem[12'hF13] = 12'hFFF;
	mem[12'hF14] = 12'hFFF;
	mem[12'hF15] = 12'hFFF;
	mem[12'hF16] = 12'hFFF;
	mem[12'hF17] = 12'hFFF;
	mem[12'hF18] = 12'hFFF;
	mem[12'hF19] = 12'hFFF;
	mem[12'hF1A] = 12'hFFF;
	mem[12'hF1B] = 12'hFFF;
	mem[12'hF1C] = 12'hFFF;
	mem[12'hF1D] = 12'hFFF;
	mem[12'hF1E] = 12'hFFF;
	mem[12'hF1F] = 12'hFFF;
	mem[12'hF20] = 12'hFFF;
	mem[12'hF21] = 12'hFFF;
	mem[12'hF22] = 12'hFFF;
	mem[12'hF23] = 12'hFFF;
	mem[12'hF24] = 12'hFFF;
	mem[12'hF25] = 12'hFFF;
	mem[12'hF26] = 12'hFFF;
	mem[12'hF27] = 12'hFFF;
	mem[12'hF28] = 12'hFFF;
	mem[12'hF29] = 12'hFFF;
	mem[12'hF2A] = 12'hFFF;
	mem[12'hF2B] = 12'hFFF;
	mem[12'hF2C] = 12'hFFF;
	mem[12'hF2D] = 12'hFFF;
	mem[12'hF2E] = 12'hFFF;
	mem[12'hF2F] = 12'hFFF;
	mem[12'hF30] = 12'hFFF;
	mem[12'hF31] = 12'hFFF;
	mem[12'hF32] = 12'hFFF;
	mem[12'hF33] = 12'hFFF;
	mem[12'hF34] = 12'hFFF;
	mem[12'hF35] = 12'hFFF;
	mem[12'hF36] = 12'hFFF;
	mem[12'hF37] = 12'hFFF;
	mem[12'hF38] = 12'hFFF;
	mem[12'hF39] = 12'hFFF;
	mem[12'hF3A] = 12'hFFF;
	mem[12'hF3B] = 12'hFFF;
	mem[12'hF3C] = 12'hFFF;
	mem[12'hF3D] = 12'hFFF;
	mem[12'hF3E] = 12'hFFF;
	mem[12'hF3F] = 12'hFFF;
	mem[12'hF40] = 12'hFFF;
	mem[12'hF41] = 12'hFFF;
	mem[12'hF42] = 12'hFFF;
	mem[12'hF43] = 12'hFFF;
	mem[12'hF44] = 12'hFFF;
	mem[12'hF45] = 12'hFFF;
	mem[12'hF46] = 12'hFFF;
	mem[12'hF47] = 12'hFFF;
	mem[12'hF48] = 12'hFFF;
	mem[12'hF49] = 12'hFFF;
	mem[12'hF4A] = 12'hFFF;
	mem[12'hF4B] = 12'hFFF;
	mem[12'hF4C] = 12'hFFF;
	mem[12'hF4D] = 12'hFFF;
	mem[12'hF4E] = 12'hFFF;
	mem[12'hF4F] = 12'hFFF;
	mem[12'hF50] = 12'hFFF;
	mem[12'hF51] = 12'hFFF;
	mem[12'hF52] = 12'hFFF;
	mem[12'hF53] = 12'hFFF;
	mem[12'hF54] = 12'hFFF;
	mem[12'hF55] = 12'hFFF;
	mem[12'hF56] = 12'hFFF;
	mem[12'hF57] = 12'hFFF;
	mem[12'hF58] = 12'hFFF;
	mem[12'hF59] = 12'hFFF;
	mem[12'hF5A] = 12'hFFF;
	mem[12'hF5B] = 12'hFFF;
	mem[12'hF5C] = 12'hFFF;
	mem[12'hF5D] = 12'hFFF;
	mem[12'hF5E] = 12'hFFF;
	mem[12'hF5F] = 12'hFFF;
	mem[12'hF60] = 12'hFFF;
	mem[12'hF61] = 12'hFFF;
	mem[12'hF62] = 12'hFFF;
	mem[12'hF63] = 12'hFFF;
	mem[12'hF64] = 12'hFFF;
	mem[12'hF65] = 12'hFFF;
	mem[12'hF66] = 12'hFFF;
	mem[12'hF67] = 12'hFFF;
	mem[12'hF68] = 12'hFFF;
	mem[12'hF69] = 12'hFFF;
	mem[12'hF6A] = 12'hFFF;
	mem[12'hF6B] = 12'hFFF;
	mem[12'hF6C] = 12'hFFF;
	mem[12'hF6D] = 12'hFFF;
	mem[12'hF6E] = 12'hFFF;
	mem[12'hF6F] = 12'hFFF;
	mem[12'hF70] = 12'hFFF;
	mem[12'hF71] = 12'hFFF;
	mem[12'hF72] = 12'hFFF;
	mem[12'hF73] = 12'hFFF;
	mem[12'hF74] = 12'hFFF;
	mem[12'hF75] = 12'hFFF;
	mem[12'hF76] = 12'hFFF;
	mem[12'hF77] = 12'hFFF;
	mem[12'hF78] = 12'hFFF;
	mem[12'hF79] = 12'hFFF;
	mem[12'hF7A] = 12'hFFF;
	mem[12'hF7B] = 12'hFFF;
	mem[12'hF7C] = 12'hFFF;
	mem[12'hF7D] = 12'hFFF;
	mem[12'hF7E] = 12'hFFF;
	mem[12'hF7F] = 12'hFFF;
	mem[12'hF80] = 12'hFFF;
	mem[12'hF81] = 12'hFFF;
	mem[12'hF82] = 12'hFFF;
	mem[12'hF83] = 12'hFFF;
	mem[12'hF84] = 12'hFFF;
	mem[12'hF85] = 12'hFFF;
	mem[12'hF86] = 12'hFFF;
	mem[12'hF87] = 12'hFFF;
	mem[12'hF88] = 12'hFFF;
	mem[12'hF89] = 12'hFFF;
	mem[12'hF8A] = 12'hFFF;
	mem[12'hF8B] = 12'hFFF;
	mem[12'hF8C] = 12'hFFF;
	mem[12'hF8D] = 12'hFFF;
	mem[12'hF8E] = 12'hFFF;
	mem[12'hF8F] = 12'hFFF;
	mem[12'hF90] = 12'hFFF;
	mem[12'hF91] = 12'hFFF;
	mem[12'hF92] = 12'hFFF;
	mem[12'hF93] = 12'hFFF;
	mem[12'hF94] = 12'hFFF;
	mem[12'hF95] = 12'hFFF;
	mem[12'hF96] = 12'hFFF;
	mem[12'hF97] = 12'hFFF;
	mem[12'hF98] = 12'hFFF;
	mem[12'hF99] = 12'hFFF;
	mem[12'hF9A] = 12'hFFF;
	mem[12'hF9B] = 12'hFFF;
	mem[12'hF9C] = 12'hFFF;
	mem[12'hF9D] = 12'hFFF;
	mem[12'hF9E] = 12'hFFF;
	mem[12'hF9F] = 12'hFFF;
	mem[12'hFA0] = 12'hFFF;
	mem[12'hFA1] = 12'hFFF;
	mem[12'hFA2] = 12'hFFF;
	mem[12'hFA3] = 12'hFFF;
	mem[12'hFA4] = 12'hFFF;
	mem[12'hFA5] = 12'hFFF;
	mem[12'hFA6] = 12'hFFF;
	mem[12'hFA7] = 12'hFFF;
	mem[12'hFA8] = 12'hFFF;
	mem[12'hFA9] = 12'hFFF;
	mem[12'hFAA] = 12'hFFF;
	mem[12'hFAB] = 12'hFFF;
	mem[12'hFAC] = 12'hFFF;
	mem[12'hFAD] = 12'hFFF;
	mem[12'hFAE] = 12'hFFF;
	mem[12'hFAF] = 12'hFFF;
	mem[12'hFB0] = 12'hFFF;
	mem[12'hFB1] = 12'hFFF;
	mem[12'hFB2] = 12'hFFF;
	mem[12'hFB3] = 12'hFFF;
	mem[12'hFB4] = 12'hFFF;
	mem[12'hFB5] = 12'hFFF;
	mem[12'hFB6] = 12'hFFF;
	mem[12'hFB7] = 12'hFFF;
	mem[12'hFB8] = 12'hFFF;
	mem[12'hFB9] = 12'hFFF;
	mem[12'hFBA] = 12'hFFF;
	mem[12'hFBB] = 12'hFFF;
	mem[12'hFBC] = 12'hFFF;
	mem[12'hFBD] = 12'hFFF;
	mem[12'hFBE] = 12'hFFF;
	mem[12'hFBF] = 12'hFFF;
	mem[12'hFC0] = 12'hFFF;
	mem[12'hFC1] = 12'hFFF;
	mem[12'hFC2] = 12'hFFF;
	mem[12'hFC3] = 12'hFFF;
	mem[12'hFC4] = 12'hFFF;
	mem[12'hFC5] = 12'hFFF;
	mem[12'hFC6] = 12'hFFF;
	mem[12'hFC7] = 12'hFFF;
	mem[12'hFC8] = 12'hFFF;
	mem[12'hFC9] = 12'hFFF;
	mem[12'hFCA] = 12'hFFF;
	mem[12'hFCB] = 12'hFFF;
	mem[12'hFCC] = 12'hFFF;
	mem[12'hFCD] = 12'hFFF;
	mem[12'hFCE] = 12'hFFF;
	mem[12'hFCF] = 12'hFFF;
	mem[12'hFD0] = 12'hFFF;
	mem[12'hFD1] = 12'hFFF;
	mem[12'hFD2] = 12'hFFF;
	mem[12'hFD3] = 12'hFFF;
	mem[12'hFD4] = 12'hFFF;
	mem[12'hFD5] = 12'hFFF;
	mem[12'hFD6] = 12'hFFF;
	mem[12'hFD7] = 12'hFFF;
	mem[12'hFD8] = 12'hFFF;
	mem[12'hFD9] = 12'hFFF;
	mem[12'hFDA] = 12'hFFF;
	mem[12'hFDB] = 12'hFFF;
	mem[12'hFDC] = 12'hFFF;
	mem[12'hFDD] = 12'hFFF;
	mem[12'hFDE] = 12'hFFF;
	mem[12'hFDF] = 12'hFFF;
	mem[12'hFE0] = 12'hFFF;
	mem[12'hFE1] = 12'hFFF;
	mem[12'hFE2] = 12'hFFF;
	mem[12'hFE3] = 12'hFFF;
	mem[12'hFE4] = 12'hFFF;
	mem[12'hFE5] = 12'hFFF;
	mem[12'hFE6] = 12'hFFF;
	mem[12'hFE7] = 12'hFFF;
	mem[12'hFE8] = 12'hFFF;
	mem[12'hFE9] = 12'hFFF;
	mem[12'hFEA] = 12'hFFF;
	mem[12'hFEB] = 12'hFFF;
	mem[12'hFEC] = 12'hFFF;
	mem[12'hFED] = 12'hFFF;
	mem[12'hFEE] = 12'hFFF;
	mem[12'hFEF] = 12'hFFF;
	mem[12'hFF0] = 12'hFFF;
	mem[12'hFF1] = 12'hFFF;
	mem[12'hFF2] = 12'hFFF;
	mem[12'hFF3] = 12'hFFF;
	mem[12'hFF4] = 12'hFFF;
	mem[12'hFF5] = 12'hFFF;
	mem[12'hFF6] = 12'hFFF;
	mem[12'hFF7] = 12'hFFF;
	mem[12'hFF8] = 12'hFFF;
	mem[12'hFF9] = 12'hFFF;
	mem[12'hFFA] = 12'hFFF;
	mem[12'hFFB] = 12'hFFF;
	mem[12'hFFC] = 12'hFFF;
	mem[12'hFFD] = 12'hFFF;
	mem[12'hFFE] = 12'hFFF;
	mem[12'hFFF] = 12'hFFF;
end

always @(posedge clock)
begin
    address_q <= address;
    q <= mem[address_q];
end
endmodule
