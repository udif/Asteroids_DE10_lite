../Drawing_priority.sv