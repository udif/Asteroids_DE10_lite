../Draw_Ghost.sv