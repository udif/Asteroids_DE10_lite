../Ghost_unit.sv