../Move_Ghost.sv